-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity trip_report is
  generic (
    INDEX_WIDTH : integer := 32;
    TAG_WIDTH   : integer := 1
  );
  port (
    kcd_clk                                       : in std_logic;
    kcd_reset                                     : in std_logic;
    input_input_valid                             : in std_logic;
    input_input_ready                             : out std_logic;
    input_input_dvalid                            : in std_logic;
    input_input_last                              : in std_logic;
    input_input                                   : in std_logic_vector(63 downto 0);
    input_input_count                             : in std_logic_vector(3 downto 0);
    input_input_unl_valid                         : in std_logic;
    input_input_unl_ready                         : out std_logic;
    input_input_unl_tag                           : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    input_input_cmd_valid                         : out std_logic;
    input_input_cmd_ready                         : in std_logic;
    input_input_cmd_firstIdx                      : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_input_cmd_lastIdx                       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_input_cmd_tag                           : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_timestamp_valid                        : out std_logic;
    output_timestamp_ready                        : in std_logic;
    output_timestamp_dvalid                       : out std_logic;
    output_timestamp_last                         : out std_logic;
    output_timestamp_length                       : out std_logic_vector(31 downto 0);
    output_timestamp_count                        : out std_logic_vector(0 downto 0);
    output_timestamp_chars_valid                  : out std_logic;
    output_timestamp_chars_ready                  : in std_logic;
    output_timestamp_chars_dvalid                 : out std_logic;
    output_timestamp_chars_last                   : out std_logic;
    output_timestamp_chars                        : out std_logic_vector(7 downto 0);
    output_timestamp_chars_count                  : out std_logic_vector(0 downto 0);
    output_timezone_valid                         : out std_logic;
    output_timezone_ready                         : in std_logic;
    output_timezone_dvalid                        : out std_logic;
    output_timezone_last                          : out std_logic;
    output_timezone                               : out std_logic_vector(63 downto 0);
    output_vin_valid                              : out std_logic;
    output_vin_ready                              : in std_logic;
    output_vin_dvalid                             : out std_logic;
    output_vin_last                               : out std_logic;
    output_vin                                    : out std_logic_vector(63 downto 0);
    output_odometer_valid                         : out std_logic;
    output_odometer_ready                         : in std_logic;
    output_odometer_dvalid                        : out std_logic;
    output_odometer_last                          : out std_logic;
    output_odometer                               : out std_logic_vector(63 downto 0);
    output_hypermiling_valid                      : out std_logic;
    output_hypermiling_ready                      : in std_logic;
    output_hypermiling_dvalid                     : out std_logic;
    output_hypermiling_last                       : out std_logic;
    output_hypermiling                            : out std_logic_vector(7 downto 0);
    output_avgspeed_valid                         : out std_logic;
    output_avgspeed_ready                         : in std_logic;
    output_avgspeed_dvalid                        : out std_logic;
    output_avgspeed_last                          : out std_logic;
    output_avgspeed                               : out std_logic_vector(63 downto 0);
    output_sec_in_band_valid                      : out std_logic;
    output_sec_in_band_ready                      : in std_logic;
    output_sec_in_band_dvalid                     : out std_logic;
    output_sec_in_band_last                       : out std_logic;
    output_sec_in_band                            : out std_logic_vector(63 downto 0);
    output_miles_in_time_range_valid              : out std_logic;
    output_miles_in_time_range_ready              : in std_logic;
    output_miles_in_time_range_dvalid             : out std_logic;
    output_miles_in_time_range_last               : out std_logic;
    output_miles_in_time_range                    : out std_logic_vector(63 downto 0);
    output_const_speed_miles_in_band_valid        : out std_logic;
    output_const_speed_miles_in_band_ready        : in std_logic;
    output_const_speed_miles_in_band_dvalid       : out std_logic;
    output_const_speed_miles_in_band_last         : out std_logic;
    output_const_speed_miles_in_band              : out std_logic_vector(63 downto 0);
    output_vary_speed_miles_in_band_valid         : out std_logic;
    output_vary_speed_miles_in_band_ready         : in std_logic;
    output_vary_speed_miles_in_band_dvalid        : out std_logic;
    output_vary_speed_miles_in_band_last          : out std_logic;
    output_vary_speed_miles_in_band               : out std_logic_vector(63 downto 0);
    output_sec_decel_valid                        : out std_logic;
    output_sec_decel_ready                        : in std_logic;
    output_sec_decel_dvalid                       : out std_logic;
    output_sec_decel_last                         : out std_logic;
    output_sec_decel                              : out std_logic_vector(63 downto 0);
    output_sec_accel_valid                        : out std_logic;
    output_sec_accel_ready                        : in std_logic;
    output_sec_accel_dvalid                       : out std_logic;
    output_sec_accel_last                         : out std_logic;
    output_sec_accel                              : out std_logic_vector(63 downto 0);
    output_braking_valid                          : out std_logic;
    output_braking_ready                          : in std_logic;
    output_braking_dvalid                         : out std_logic;
    output_braking_last                           : out std_logic;
    output_braking                                : out std_logic_vector(63 downto 0);
    output_accel_valid                            : out std_logic;
    output_accel_ready                            : in std_logic;
    output_accel_dvalid                           : out std_logic;
    output_accel_last                             : out std_logic;
    output_accel                                  : out std_logic_vector(63 downto 0);
    output_orientation_valid                      : out std_logic;
    output_orientation_ready                      : in std_logic;
    output_orientation_dvalid                     : out std_logic;
    output_orientation_last                       : out std_logic;
    output_orientation                            : out std_logic_vector(7 downto 0);
    output_small_speed_var_valid                  : out std_logic;
    output_small_speed_var_ready                  : in std_logic;
    output_small_speed_var_dvalid                 : out std_logic;
    output_small_speed_var_last                   : out std_logic;
    output_small_speed_var                        : out std_logic_vector(63 downto 0);
    output_large_speed_var_valid                  : out std_logic;
    output_large_speed_var_ready                  : in std_logic;
    output_large_speed_var_dvalid                 : out std_logic;
    output_large_speed_var_last                   : out std_logic;
    output_large_speed_var                        : out std_logic_vector(63 downto 0);
    output_accel_decel_valid                      : out std_logic;
    output_accel_decel_ready                      : in std_logic;
    output_accel_decel_dvalid                     : out std_logic;
    output_accel_decel_last                       : out std_logic;
    output_accel_decel                            : out std_logic_vector(63 downto 0);
    output_speed_changes_valid                    : out std_logic;
    output_speed_changes_ready                    : in std_logic;
    output_speed_changes_dvalid                   : out std_logic;
    output_speed_changes_last                     : out std_logic;
    output_speed_changes                          : out std_logic_vector(63 downto 0);
    output_timestamp_unl_valid                    : in std_logic;
    output_timestamp_unl_ready                    : out std_logic;
    output_timestamp_unl_tag                      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_timezone_unl_valid                     : in std_logic;
    output_timezone_unl_ready                     : out std_logic;
    output_timezone_unl_tag                       : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_vin_unl_valid                          : in std_logic;
    output_vin_unl_ready                          : out std_logic;
    output_vin_unl_tag                            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_odometer_unl_valid                     : in std_logic;
    output_odometer_unl_ready                     : out std_logic;
    output_odometer_unl_tag                       : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_hypermiling_unl_valid                  : in std_logic;
    output_hypermiling_unl_ready                  : out std_logic;
    output_hypermiling_unl_tag                    : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_avgspeed_unl_valid                     : in std_logic;
    output_avgspeed_unl_ready                     : out std_logic;
    output_avgspeed_unl_tag                       : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_sec_in_band_unl_valid                  : in std_logic;
    output_sec_in_band_unl_ready                  : out std_logic;
    output_sec_in_band_unl_tag                    : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_miles_in_time_range_unl_valid          : in std_logic;
    output_miles_in_time_range_unl_ready          : out std_logic;
    output_miles_in_time_range_unl_tag            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_const_speed_miles_in_band_unl_valid    : in std_logic;
    output_const_speed_miles_in_band_unl_ready    : out std_logic;
    output_const_speed_miles_in_band_unl_tag      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_vary_speed_miles_in_band_unl_valid     : in std_logic;
    output_vary_speed_miles_in_band_unl_ready     : out std_logic;
    output_vary_speed_miles_in_band_unl_tag       : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_sec_decel_unl_valid                    : in std_logic;
    output_sec_decel_unl_ready                    : out std_logic;
    output_sec_decel_unl_tag                      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_sec_accel_unl_valid                    : in std_logic;
    output_sec_accel_unl_ready                    : out std_logic;
    output_sec_accel_unl_tag                      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_braking_unl_valid                      : in std_logic;
    output_braking_unl_ready                      : out std_logic;
    output_braking_unl_tag                        : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_accel_unl_valid                        : in std_logic;
    output_accel_unl_ready                        : out std_logic;
    output_accel_unl_tag                          : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_orientation_unl_valid                  : in std_logic;
    output_orientation_unl_ready                  : out std_logic;
    output_orientation_unl_tag                    : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_small_speed_var_unl_valid              : in std_logic;
    output_small_speed_var_unl_ready              : out std_logic;
    output_small_speed_var_unl_tag                : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_large_speed_var_unl_valid              : in std_logic;
    output_large_speed_var_unl_ready              : out std_logic;
    output_large_speed_var_unl_tag                : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_accel_decel_unl_valid                  : in std_logic;
    output_accel_decel_unl_ready                  : out std_logic;
    output_accel_decel_unl_tag                    : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_speed_changes_unl_valid                : in std_logic;
    output_speed_changes_unl_ready                : out std_logic;
    output_speed_changes_unl_tag                  : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_timestamp_cmd_valid                    : out std_logic;
    output_timestamp_cmd_ready                    : in std_logic;
    output_timestamp_cmd_firstIdx                 : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_timestamp_cmd_lastIdx                  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_timestamp_cmd_tag                      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_timezone_cmd_valid                     : out std_logic;
    output_timezone_cmd_ready                     : in std_logic;
    output_timezone_cmd_firstIdx                  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_timezone_cmd_lastIdx                   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_timezone_cmd_tag                       : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_vin_cmd_valid                          : out std_logic;
    output_vin_cmd_ready                          : in std_logic;
    output_vin_cmd_firstIdx                       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_vin_cmd_lastIdx                        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_vin_cmd_tag                            : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_odometer_cmd_valid                     : out std_logic;
    output_odometer_cmd_ready                     : in std_logic;
    output_odometer_cmd_firstIdx                  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_odometer_cmd_lastIdx                   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_odometer_cmd_tag                       : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_hypermiling_cmd_valid                  : out std_logic;
    output_hypermiling_cmd_ready                  : in std_logic;
    output_hypermiling_cmd_firstIdx               : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_hypermiling_cmd_lastIdx                : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_hypermiling_cmd_tag                    : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_avgspeed_cmd_valid                     : out std_logic;
    output_avgspeed_cmd_ready                     : in std_logic;
    output_avgspeed_cmd_firstIdx                  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_avgspeed_cmd_lastIdx                   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_avgspeed_cmd_tag                       : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_sec_in_band_cmd_valid                  : out std_logic;
    output_sec_in_band_cmd_ready                  : in std_logic;
    output_sec_in_band_cmd_firstIdx               : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_sec_in_band_cmd_lastIdx                : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_sec_in_band_cmd_tag                    : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_miles_in_time_range_cmd_valid          : out std_logic;
    output_miles_in_time_range_cmd_ready          : in std_logic;
    output_miles_in_time_range_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_miles_in_time_range_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_miles_in_time_range_cmd_tag            : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_const_speed_miles_in_band_cmd_valid    : out std_logic;
    output_const_speed_miles_in_band_cmd_ready    : in std_logic;
    output_const_speed_miles_in_band_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_const_speed_miles_in_band_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_const_speed_miles_in_band_cmd_tag      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_vary_speed_miles_in_band_cmd_valid     : out std_logic;
    output_vary_speed_miles_in_band_cmd_ready     : in std_logic;
    output_vary_speed_miles_in_band_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_vary_speed_miles_in_band_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_vary_speed_miles_in_band_cmd_tag       : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_sec_decel_cmd_valid                    : out std_logic;
    output_sec_decel_cmd_ready                    : in std_logic;
    output_sec_decel_cmd_firstIdx                 : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_sec_decel_cmd_lastIdx                  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_sec_decel_cmd_tag                      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_sec_accel_cmd_valid                    : out std_logic;
    output_sec_accel_cmd_ready                    : in std_logic;
    output_sec_accel_cmd_firstIdx                 : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_sec_accel_cmd_lastIdx                  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_sec_accel_cmd_tag                      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_braking_cmd_valid                      : out std_logic;
    output_braking_cmd_ready                      : in std_logic;
    output_braking_cmd_firstIdx                   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_braking_cmd_lastIdx                    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_braking_cmd_tag                        : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_accel_cmd_valid                        : out std_logic;
    output_accel_cmd_ready                        : in std_logic;
    output_accel_cmd_firstIdx                     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_accel_cmd_lastIdx                      : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_accel_cmd_tag                          : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_orientation_cmd_valid                  : out std_logic;
    output_orientation_cmd_ready                  : in std_logic;
    output_orientation_cmd_firstIdx               : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_orientation_cmd_lastIdx                : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_orientation_cmd_tag                    : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_small_speed_var_cmd_valid              : out std_logic;
    output_small_speed_var_cmd_ready              : in std_logic;
    output_small_speed_var_cmd_firstIdx           : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_small_speed_var_cmd_lastIdx            : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_small_speed_var_cmd_tag                : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_large_speed_var_cmd_valid              : out std_logic;
    output_large_speed_var_cmd_ready              : in std_logic;
    output_large_speed_var_cmd_firstIdx           : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_large_speed_var_cmd_lastIdx            : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_large_speed_var_cmd_tag                : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_accel_decel_cmd_valid                  : out std_logic;
    output_accel_decel_cmd_ready                  : in std_logic;
    output_accel_decel_cmd_firstIdx               : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_accel_decel_cmd_lastIdx                : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_accel_decel_cmd_tag                    : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_speed_changes_cmd_valid                : out std_logic;
    output_speed_changes_cmd_ready                : in std_logic;
    output_speed_changes_cmd_firstIdx             : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_speed_changes_cmd_lastIdx              : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_speed_changes_cmd_tag                  : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    start                                         : in std_logic;
    stop                                          : in std_logic;
    reset                                         : in std_logic;
    idle                                          : out std_logic;
    busy                                          : out std_logic;
    done                                          : out std_logic;
    result                                        : out std_logic_vector(63 downto 0);
    input_firstidx                                : in std_logic_vector(31 downto 0);
    input_lastidx                                 : in std_logic_vector(31 downto 0);
    output_firstidx                               : in std_logic_vector(31 downto 0);
    output_lastidx                                : in std_logic_vector(31 downto 0);
    ext_platform_complete_req                     : out std_logic;
    ext_platform_complete_ack                     : in std_logic
  );
end entity;

architecture Implementation of trip_report is
begin

  battery_status_parser : BattSchemaParser
  generic map(
    EPC                                    => 8,

    -- 
    -- INTEGER FIELDS
    --
    TIMEZONE_INT_WIDTH                     => 16,
    TIMEZONE_INT_P_PIPELINE_STAGES         => 1,
    TIMEZONE_BUFFER_D                      => 1,

    VIN_INT_WIDTH                          => 16,
    VIN_INT_P_PIPELINE_STAGES              => 1,
    VIN_BUFFER_D                           => 1,

    ODOMETER_INT_WIDTH                     => 16,
    ODOMETER_INT_P_PIPELINE_STAGES         => 1,
    ODOMETER_BUFFER_D                      => 1,

    AVG_SPEED_INT_WIDTH                    => 16,
    AVG_SPEED_INT_P_PIPELINE_STAGES        => 1,
    AVG_SPEED_BUFFER_D                     => 1,

    S_ACC_DEC_INT_WIDTH                    => 16,
    S_ACC_DEC_INT_P_PIPELINE_STAGES        => 1,
    S_ACC_DEC_BUFFER_D                     => 1,

    E_SPD_CHG_INT_WIDTH                    => 16,
    E_SPD_CHG_INT_P_PIPELINE_STAGES        => 1,
    E_SPD_CHG_BUFFER_D                     => 1,

    -- 
    -- BOOLEAN FIELDS
    --
    HYPER_MILING_BUFFER_D                  => 1,
    ORIENTATION_BUFFER_D                   => 1,

    -- 
    -- INTEGER ARRAY FIELDS
    --
    SECS_IN_B_INT_WIDTH                    => 16,
    SECS_IN_B_INT_P_PIPELINE_STAGES        => 1,
    SECS_IN_B_BUFFER_D                     => 1,

    MILES_IN_TIME_INT_WIDTH                => 16,
    MILES_IN_TIME_INT_P_PIPELINE_STAGES    => 1,
    MILES_IN_TIME_BUFFER_D                 => 1,
    CONST_SPD_M_IN_B_INT_WIDTH             => 16,
    CONST_SPD_M_IN_B_INT_P_PIPELINE_STAGES => 1,
    CONST_SPD_M_IN_B_BUFFER_D              => 1,
    VAR_SPD_M_IN_B_INT_WIDTH               => 16,
    VAR_SPD_M_IN_B_INT_P_PIPELINE_STAGES   => 1,
    VAR_SPD_M_IN_B_BUFFER_D                => 1,
    SECONDS_DECEL_INT_WIDTH                => 16,
    SECONDS_DECEL_INT_P_PIPELINE_STAGES    => 1,
    SECONDS_DECEL_BUFFER_D                 => 1,
    SECONDS_ACCEL_INT_WIDTH                => 16,
    SECONDS_ACCEL_INT_P_PIPELINE_STAGES    => 1,
    SECONDS_ACCEL_BUFFER_D                 => 1,
    BRK_M_T_10S_INT_WIDTH                  => 16,
    BRK_M_T_10S_INT_P_PIPELINE_STAGES      => 1,
    BRK_M_T_10S_BUFFER_D                   => 1,
    ACCEL_M_T_10S_INT_WIDTH                => 16,
    ACCEL_M_T_10S_INT_P_PIPELINE_STAGES    => 1,
    ACCEL_M_T_10S_BUFFER_D                 => 1,
    SMALL_SPD_V_M_INT_WIDTH                => 16,
    SMALL_SPD_V_M_INT_P_PIPELINE_STAGES    => 1,
    SMALL_SPD_V_M_BUFFER_D                 => 1,
    LARGE_SPD_V_M_INT_WIDTH                => 16,
    LARGE_SPD_V_M_INT_P_PIPELINE_STAGES    => 1,
    LARGE_SPD_V_M_BUFFER_D                 => 1,

    -- 
    -- STRING FIELDS
    --
    TIMESTAMP_BUFFER_D                     => 1,

    END_REQ_EN                             => false
  );
  port map(
    clk                    => open,
    reset                  => open,

    in_valid               => open,
    in_ready               => open,
    in_data                => open,
    in_last                => open,
    in_stai                => open,
    in_endi                => open,
    in_strb                => open,

    end_req                => open,
    end_ack                => open,

    timezone_valid         => open,
    timezone_ready         => open,
    timezone_data          => open,
    timezone_strb          => open,
    timezone_last          => open,

    --    
    -- INTEGER FIELDS   
    --    
    vin_valid              => open,
    vin_ready              => open,
    vin_data               => open,
    vin_strb               => open,
    vin_last               => open,

    odometer_valid         => open,
    odometer_ready         => open,
    odometer_data          => open,
    odometer_strb          => open,
    odometer_last          => open,

    avg_speed_valid        => open,
    avg_speed_ready        => open,
    avg_speed_data         => open,
    avg_speed_strb         => open,
    avg_speed_last         => open,

    s_acc_dec_valid        => open,
    s_acc_dec_ready        => open,
    s_acc_dec_data         => open,
    s_acc_dec_strb         => open,
    s_acc_dec_last         => open,

    e_spd_chg_valid        => open,
    e_spd_chg_ready        => open,
    e_spd_chg_data         => open,
    e_spd_chg_strb         => open,
    e_spd_chg_last         => open,

    --    
    -- BOOLEAN FIELDS   
    --    
    hyper_miling_valid     => open,
    hyper_miling_ready     => open,
    hyper_miling_data      => open,
    hyper_miling_strb      => open,
    hyper_miling_last      => open,

    orientation_valid      => open,
    orientation_ready      => open,
    orientation_data       => open,
    orientation_strb       => open,
    orientation_last       => open,

    --    
    -- INTEGER ARRAY FIELDS   
    --    
    secs_in_b_valid        => open,
    secs_in_b_ready        => open,
    secs_in_b_data         => open,
    secs_in_b_strb         => open,
    secs_in_b_last         => open,

    miles_in_time_valid    => open,
    miles_in_time_ready    => open,
    miles_in_time_data     => open,
    miles_in_time_strb     => open,
    miles_in_time_last     => open,
    const_spd_m_in_b_valid => open,
    const_spd_m_in_b_ready => open,
    const_spd_m_in_b_data  => open,
    const_spd_m_in_b_strb  => open,
    const_spd_m_in_b_last  => open,
    var_spd_m_in_b_valid   => open,
    var_spd_m_in_b_ready   => open,
    var_spd_m_in_b_data    => open,
    var_spd_m_in_b_strb    => open,
    var_spd_m_in_b_last    => open,
    seconds_decel_valid    => open,
    seconds_decel_ready    => open,
    seconds_decel_data     => open,
    seconds_decel_strb     => open,
    seconds_decel_last     => open,
    seconds_accel_valid    => open,
    seconds_accel_ready    => open,
    seconds_accel_data     => open,
    seconds_accel_strb     => open,
    seconds_accel_last     => open,
    brk_m_t_10s_valid      => open,
    brk_m_t_10s_ready      => open,
    brk_m_t_10s_data       => open,
    brk_m_t_10s_strb       => open,
    brk_m_t_10s_last       => open,
    accel_m_t_10s_valid    => open,
    accel_m_t_10s_ready    => open,
    accel_m_t_10s_data     => open,
    accel_m_t_10s_strb     => open,
    accel_m_t_10s_last     => open,
    small_spd_v_m_valid    => open,
    small_spd_v_m_ready    => open,
    small_spd_v_m_data     => open,
    small_spd_v_m_strb     => open,
    small_spd_v_m_last     => open,
    large_spd_v_m_valid    => open,
    large_spd_v_m_ready    => open,
    large_spd_v_m_data     => open,
    large_spd_v_m_strb     => open,
    large_spd_v_m_last     => open,

    --    
    -- STRING FIELDS   
    -- 
    timestamp_valid        => open,
    timestamp_ready        => open,
    timestamp_data         => open,
    timestamp_last         => open,
    timestamp_stai         => open,
    timestamp_endi         => open,
    timestamp_strb         => open
  );

end architecture;