-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.battery_status_pkg.all;
use work.Stream_pkg.all;

entity battery_status_sub is
  generic (
    INDEX_WIDTH : integer := 32;
    TAG_WIDTH   : integer := 1
  );
  port (
    kcd_clk                     : in std_logic;
    kcd_reset                   : in std_logic;
    input_input_valid           : in std_logic;
    input_input_ready           : out std_logic;
    input_input_dvalid          : in std_logic;
    input_input_last            : in std_logic;
    input_input                 : in std_logic_vector(63 downto 0);
    input_input_count           : in std_logic_vector(3 downto 0);
    input_input_unl_valid       : in std_logic;
    input_input_unl_ready       : out std_logic;
    input_input_unl_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    input_input_cmd_valid       : out std_logic;
    input_input_cmd_ready       : in std_logic;
    input_input_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_input_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_input_cmd_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_voltage_valid        : out std_logic;
    output_voltage_ready        : in std_logic;
    output_voltage_dvalid       : out std_logic;
    output_voltage_last         : out std_logic;
    output_voltage_length       : out std_logic_vector(31 downto 0);
    output_voltage_count        : out std_logic_vector(0 downto 0);
    output_voltage_item_valid   : out std_logic;
    output_voltage_item_ready   : in std_logic;
    output_voltage_item_dvalid  : out std_logic;
    output_voltage_item_last    : out std_logic;
    output_voltage_item         : out std_logic_vector(63 downto 0);
    output_voltage_item_count   : out std_logic_vector(0 downto 0);
    output_voltage_unl_valid    : in std_logic;
    output_voltage_unl_ready    : out std_logic;
    output_voltage_unl_tag      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_voltage_cmd_valid    : out std_logic;
    output_voltage_cmd_ready    : in std_logic;
    output_voltage_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_voltage_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_voltage_cmd_tag      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    start                       : in std_logic;
    stop                        : in std_logic;
    reset                       : in std_logic;
    idle                        : out std_logic;
    busy                        : out std_logic;
    done                        : out std_logic;
    result                      : out std_logic_vector(63 downto 0);
    input_firstidx              : in std_logic_vector(31 downto 0);
    input_lastidx               : in std_logic_vector(31 downto 0);
    output_firstidx             : in std_logic_vector(31 downto 0);
    output_lastidx              : in std_logic_vector(31 downto 0)
  );
end entity;

architecture Implementation of battery_status_sub is

  -- elements per cycle of input stream
  -- matches the value set in the schema (generate.py)
  constant EPC : natural := 8;

  type state_t is (
    STATE_IDLE,         -- idle
    STATE_REQ_READ,     -- send read request
    STATE_REQ_WRITE,    -- send write request
    STATE_UNLOCK_READ,  -- unlock read
    STATE_UNLOCK_WRITE, -- unlock write
    STATE_DONE          -- done
  );

  -- state signals
  signal state, state_next     : state_t;

  -- parser output signals
  signal json_out_valid        : std_logic;
  signal json_out_ready        : std_logic;
  signal json_out_data         : std_logic_vector(63 downto 0);
  signal json_out_last         : std_logic_vector(2 downto 0);
  signal json_out_strb         : std_logic;

  signal int_input_input_ready : std_logic;

  signal strb                  : std_logic_vector(EPC - 1 downto 0);
  signal int_in_last           : std_logic_vector(2 * EPC - 1 downto 0);

  signal cmd_complete          : std_logic;

  signal record_counter        : unsigned(63 downto 0);

begin

  counter : process (kcd_clk)
    is
  begin
    if rising_edge(kcd_clk) then
      if json_out_ready = '1' and json_out_valid = '1' and json_out_last(1) = '1' then
        record_counter <= record_counter + 1;
      end if;
      if kcd_reset = '1' or reset = '1' then
        record_counter <= (others => '0');
      end if;
    end if;
  end process;

  result <= std_logic_vector(record_counter);

  comb : process (
    start,
    reset,
    state,
    input_firstidx,
    input_lastidx,
    output_firstidx,
    output_lastidx,
    int_input_input_ready,
    input_input_cmd_ready,
    output_voltage_cmd_ready,
    input_input_unl_valid,
    output_voltage_unl_valid
    ) is
  begin

    -- read request defaults
    input_input_cmd_valid       <= '0';
    input_input_cmd_firstIdx    <= input_firstidx;
    input_input_cmd_lastIdx     <= input_lastidx;
    input_input_cmd_tag         <= (others => '0');
    input_input_unl_ready       <= '0';

    -- write request defaults
    output_voltage_cmd_valid    <= '0';
    output_voltage_cmd_firstIdx <= output_firstidx;
    output_voltage_cmd_lastIdx  <= output_lastidx;
    output_voltage_cmd_tag      <= (others => '0');
    output_voltage_unl_ready    <= '0';

    -- next state is the same if not changed
    state_next                  <= state;

    -- internal signal
    input_input_ready           <= int_input_input_ready;

    case state is

        -- wait for start signal
      when STATE_IDLE =>
        done <= '0';
        busy <= '0';
        idle <= '1';

        if start = '1' then
          state_next <= STATE_REQ_READ;
        end if;

        -- send read request
      when STATE_REQ_READ =>
        done                  <= '0';
        busy                  <= '1';
        idle                  <= '0';

        input_input_cmd_valid <= '1';

        -- handshake
        if input_input_cmd_ready = '1' then
          state_next <= STATE_REQ_WRITE;
        end if;

        -- send write request
      when STATE_REQ_WRITE =>
        done                     <= '0';
        busy                     <= '1';
        idle                     <= '0';

        output_voltage_cmd_valid <= '1';

        -- handshake
        if output_voltage_cmd_ready = '1' then
          state_next <= STATE_UNLOCK_READ;
        end if;

        -- unlock read
      when STATE_UNLOCK_READ =>
        done <= '0';
        busy <= '1';
        idle <= '0';

        if input_input_unl_valid = '1' then
          input_input_unl_ready <= '1';
          state_next            <= STATE_UNLOCK_WRITE;
        end if;

        -- unlock write
      when STATE_UNLOCK_WRITE =>
        done <= '0';
        busy <= '1';
        idle <= '0';

        if output_voltage_unl_valid = '1' then
          output_voltage_unl_ready <= '1';
          state_next               <= STATE_DONE;
        end if;

        -- wait for kernel reset
      when STATE_DONE =>
        done <= '1';
        busy <= '0';
        idle <= '1';

        if reset = '1' then
          state_next <= STATE_IDLE;
        end if;

    end case;

  end process;

  seq : process (kcd_clk)
  begin
    if rising_edge(kcd_clk) then
      state <= state_next;

      if kcd_reset = '1' then
        state <= STATE_IDLE;
      end if;

    end if;
  end process;

  tydi_strb : process (input_input_dvalid, input_input_count)
  begin
    strb <= (others => '0');
    for i in strb'range loop
      if unsigned(input_input_count) = 0 or i < unsigned(input_input_count) then
        strb(i) <= input_input_dvalid;
      end if;
    end loop;
  end process;

  int_in_last_proc : process (input_input_last)
  begin
    int_in_last              <= (others => '0');
    -- all records are currently sent in one transfer, so there's no difference
    -- between the two dimensions going into the parser.
    int_in_last(EPC * 2 - 2) <= input_input_last;
    int_in_last(EPC * 2 - 1) <= input_input_last;
  end process;

  battery_status_parser : BattSchemaParser
  generic map(
    EPC                   => EPC,
    INT_WIDTH             => 64,
    INT_P_PIPELINE_STAGES => 4,
    END_REQ_EN            => false
  )
  port map(
    clk       => kcd_clk,
    reset     => kcd_reset,
    in_valid  => input_input_valid,
    in_ready  => int_input_input_ready,
    in_data   => input_input,
    in_last   => int_in_last,
    in_stai => (others => '0'),
    in_endi => (others => '1'),
    in_strb   => strb,
    end_req   => '0',  -- not implemented
    end_ack   => open, -- not implemented
    out_valid => json_out_valid,
    out_ready => json_out_ready,
    out_data  => json_out_data,
    out_last  => json_out_last,
    out_strb  => json_out_strb
  );

  convert_proc : process (kcd_clk) is

    type input_holding_reg_type is record
      valid         : std_logic;
      dvalid        : std_logic;
      data          : std_logic_vector(63 downto 0);
      end_of_array  : std_logic;
      end_of_object : std_logic;
      end_of_query  : std_logic;
    end record;
    variable i : input_holding_reg_type;

    type count_output_holding_reg_type is record
      valid  : std_logic;
      dvalid : std_logic;
      data   : std_logic_vector(31 downto 0);
      last   : std_logic;
    end record;
    variable oc : count_output_holding_reg_type;

    type element_output_holding_reg_type is record
      valid  : std_logic;
      dvalid : std_logic;
      data   : std_logic_vector(63 downto 0);
      last   : std_logic;
    end record;
    variable oe    : element_output_holding_reg_type;

    -- Current element count for length stream.
    variable count : unsigned(31 downto 0) := (others => '0');

  begin
    if rising_edge(kcd_clk) then
      cmd_complete <= '0';

      if i.valid = '0' then
        i.valid         := json_out_valid;
        i.dvalid        := json_out_strb;
        i.data          := json_out_data;
        i.end_of_array  := json_out_last(0);
        i.end_of_object := json_out_last(1);
        i.end_of_query  := json_out_last(2);
      end if;

      if output_voltage_ready = '1' then
        oc.valid := '0';
      end if;

      if output_voltage_item_ready = '1' then
        oe.valid := '0';
      end if;

      if i.valid = '1' and oc.valid = '0' and oe.valid = '0' then
        oe.dvalid := '0';
        oe.last   := '0';
        oc.dvalid := '0';
        oc.last   := '0';

        -- If the data is valid, forward it and increment the element counter.
        if i.dvalid = '1' then
          -- oe.valid  := '1';
          oe.dvalid := '1';
          oe.data   := i.data;
          count     := count + 1;
        end if;

        -- If this is the end of the current JSON object, send last to the
        -- element stream and send the element count to the length stream.
        -- We could also use end_of_array here; for valid JSON these should be
        -- equivalent.
        if i.end_of_object = '1' then
          -- oc.valid  := '1';
          oc.dvalid := '1';
          oc.data   := std_logic_vector(count);
          count     := (others => '0');
        end if;

        -- If this is the end of the current command, send last to the length
        -- stream, and send a strobe to the state machine that indicates
        -- completion.
        if i.end_of_query = '1' then
          -- oe.valid := '1';
          oe.last := '1';
          -- oc.valid := '1';
          oc.last := '1';
          cmd_complete <= '1';
        end if;

        oe.valid := i.dvalid or i.end_of_query;
        oc.valid := i.end_of_object or i.end_of_query;

        -- clear holding register
        i.valid  := '0';

      end if;

      if kcd_reset = '1' then
        i.valid  := '0';
        oc.valid := '0';
        oe.valid := '0';
        count    := (others => '0');
        cmd_complete <= '0';
      end if;

      json_out_ready             <= not i.valid;

      output_voltage_valid       <= oc.valid;
      output_voltage_dvalid      <= oc.dvalid;
      output_voltage_last        <= oc.last;
      output_voltage_length      <= oc.data;
      output_voltage_count       <= "1";

      output_voltage_item_valid  <= oe.valid;
      output_voltage_item_dvalid <= oe.dvalid;
      output_voltage_item_last   <= oe.last;
      output_voltage_item        <= oe.data;
      output_voltage_item_count  <= "1";

    end if;
  end process;

end architecture;