-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity primmap is
  generic (
    INDEX_WIDTH : integer := 32;
    TAG_WIDTH   : integer := 1
  );
  port (
    kcd_clk                 : in  std_logic;
    kcd_reset               : in  std_logic;
    in_number_valid         : in  std_logic;
    in_number_ready         : out std_logic;
    in_number_dvalid        : in  std_logic;
    in_number_last          : in  std_logic;
    in_number               : in  std_logic_vector(63 downto 0);
    in_number_unl_valid     : in  std_logic;
    in_number_unl_ready     : out std_logic;
    in_number_unl_tag       : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    in_number_cmd_valid     : out std_logic;
    in_number_cmd_ready     : in  std_logic;
    in_number_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    in_number_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    in_number_cmd_tag       : out std_logic_vector(TAG_WIDTH-1 downto 0);
    out_number_valid        : out std_logic;
    out_number_ready        : in  std_logic;
    out_number_dvalid       : out std_logic;
    out_number_last         : out std_logic;
    out_number              : out std_logic_vector(63 downto 0);
    out_number_unl_valid    : in  std_logic;
    out_number_unl_ready    : out std_logic;
    out_number_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    out_number_cmd_valid    : out std_logic;
    out_number_cmd_ready    : in  std_logic;
    out_number_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    out_number_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    out_number_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    start                   : in  std_logic;
    stop                    : in  std_logic;
    reset                   : in  std_logic;
    idle                    : out std_logic;
    busy                    : out std_logic;
    done                    : out std_logic;
    result                  : out std_logic_vector(63 downto 0);
    in_firstidx             : in  std_logic_vector(31 downto 0);
    in_lastidx              : in  std_logic_vector(31 downto 0);
    out_firstidx            : in  std_logic_vector(31 downto 0);
    out_lastidx             : in  std_logic_vector(31 downto 0)
  );
end entity;

architecture Implementation of PrimMap is
  type state_t is (STATE_IDLE,
    STATE_COMMAND_IN,
    STATE_COMMAND_OUT,
    STATE_STREAMING,
    STATE_UNLOCK_IN,
    STATE_UNLOCK_OUT,
    STATE_PLATFORM,
    STATE_DONE);

  signal state, state_next : state_t;
begin
  combinatorial_proc : process (
    in_number,
    in_number_last,
    in_number_dvalid,
    state,
    start,
    in_firstIdx,
    in_lastIdx,
    in_number_cmd_ready,
    out_firstIdx,
    out_lastIdx,
    out_number_cmd_ready,
    out_number_ready,
    in_number_valid,
    in_number_unl_valid,
    out_number_unl_valid,
    ext_platform_complete_ack,
    reset
    ) is
  begin
    in_number_cmd_valid       <= '0';
    in_number_cmd_firstIdx    <= (others => '0');
    in_number_cmd_lastIdx     <= (others => '0');
    in_number_cmd_tag         <= (others => '0');

    in_number_unl_ready       <= '0';

    in_number_ready           <= '0';

    out_number_cmd_valid      <= '0';
    out_number_cmd_firstIdx   <= (others => '0');
    out_number_cmd_lastIdx    <= (others => '0');
    out_number_cmd_tag        <= (others => '0');

    out_number_unl_ready      <= '0';

    out_number_valid          <= '0';
    out_number                <= std_logic_vector(unsigned(in_number) + 1);
    out_number_last           <= in_number_last;
    out_number_dvalid         <= in_number_dvalid;

    state_next                <= state;

    case state is
      when STATE_IDLE =>
        done <= '0';
        busy <= '0';
        idle <= '1';

        if start = '1' then
          state_next <= STATE_COMMAND_IN;
        end if;

      when STATE_COMMAND_IN =>
        done                   <= '0';
        busy                   <= '1';
        idle                   <= '0';

        in_number_cmd_valid    <= '1';
        in_number_cmd_firstIdx <= in_firstIdx;
        in_number_cmd_lastIdx  <= in_lastIdx;
        in_number_cmd_tag      <= (others => '0');

        if in_number_cmd_ready = '1' then
          state_next <= STATE_COMMAND_OUT;
        end if;

      when STATE_COMMAND_OUT =>
        done                    <= '0';
        busy                    <= '1';
        idle                    <= '0';

        out_number_cmd_valid    <= '1';
        out_number_cmd_firstIdx <= out_firstIdx;
        out_number_cmd_lastIdx  <= out_lastIdx;
        out_number_cmd_tag      <= (others => '0');

        if out_number_cmd_ready = '1' then
          state_next <= STATE_STREAMING;
        end if;

      when STATE_STREAMING =>
        done             <= '0';
        busy             <= '1';
        idle             <= '0';

        in_number_ready  <= out_number_ready;
        out_number_valid <= in_number_valid;

        -- Wait for last handshake.
        if in_number_valid = '1' and
          in_number_last = '1' and
          out_number_ready = '1'
          then
          state_next <= STATE_UNLOCK_IN;
        end if;

      when STATE_UNLOCK_IN =>
        done                <= '0';
        busy                <= '1';
        idle                <= '0';

        in_number_unl_ready <= '1';
        if in_number_unl_valid = '1' then
          state_next <= STATE_UNLOCK_OUT;
        end if;

      when STATE_UNLOCK_OUT =>
        done                 <= '0';
        busy                 <= '1';
        idle                 <= '0';

        out_number_unl_ready <= '1';
        if out_number_unl_valid = '1' then
          state_next <= STATE_PLATFORM;
        end if;

      when STATE_DONE =>
        done <= '1';
        busy <= '0';
        idle <= '1';

        if reset = '1' then
          state_next <= STATE_IDLE;
        end if;

    end case;
  end process;
  -- Sequential part:
  sequential_proc : process (kcd_clk)
  begin
    if rising_edge(kcd_clk) then
      state <= state_next;

      if kcd_reset = '1' then
        state <= STATE_IDLE;
      end if;
    end if;
  end process;
end architecture;
