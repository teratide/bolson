-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;

entity battery_status_output is
  generic (
    INDEX_WIDTH                       : integer := 32;
    TAG_WIDTH                         : integer := 1;
    OUTPUT_VOLTAGE_BUS_ADDR_WIDTH     : integer := 64;
    OUTPUT_VOLTAGE_BUS_DATA_WIDTH     : integer := 512;
    OUTPUT_VOLTAGE_BUS_LEN_WIDTH      : integer := 8;
    OUTPUT_VOLTAGE_BUS_BURST_STEP_LEN : integer := 1;
    OUTPUT_VOLTAGE_BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk                        : in std_logic;
    bcd_reset                      : in std_logic;
    kcd_clk                        : in std_logic;
    kcd_reset                      : in std_logic;
    output_voltage_valid           : in std_logic;
    output_voltage_ready           : out std_logic;
    output_voltage_dvalid          : in std_logic;
    output_voltage_last            : in std_logic;
    output_voltage_length          : in std_logic_vector(31 downto 0);
    output_voltage_count           : in std_logic_vector(0 downto 0);
    output_voltage_item_valid      : in std_logic;
    output_voltage_item_ready      : out std_logic;
    output_voltage_item_dvalid     : in std_logic;
    output_voltage_item_last       : in std_logic;
    output_voltage_item            : in std_logic_vector(63 downto 0);
    output_voltage_item_count      : in std_logic_vector(0 downto 0);
    output_voltage_bus_wreq_valid  : out std_logic;
    output_voltage_bus_wreq_ready  : in std_logic;
    output_voltage_bus_wreq_addr   : out std_logic_vector(OUTPUT_VOLTAGE_BUS_ADDR_WIDTH - 1 downto 0);
    output_voltage_bus_wreq_len    : out std_logic_vector(OUTPUT_VOLTAGE_BUS_LEN_WIDTH - 1 downto 0);
    output_voltage_bus_wdat_valid  : out std_logic;
    output_voltage_bus_wdat_ready  : in std_logic;
    output_voltage_bus_wdat_data   : out std_logic_vector(OUTPUT_VOLTAGE_BUS_DATA_WIDTH - 1 downto 0);
    output_voltage_bus_wdat_strobe : out std_logic_vector(OUTPUT_VOLTAGE_BUS_DATA_WIDTH/8 - 1 downto 0);
    output_voltage_bus_wdat_last   : out std_logic;
    output_voltage_cmd_valid       : in std_logic;
    output_voltage_cmd_ready       : out std_logic;
    output_voltage_cmd_firstIdx    : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_voltage_cmd_lastIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_voltage_cmd_ctrl        : in std_logic_vector(OUTPUT_VOLTAGE_BUS_ADDR_WIDTH * 2 - 1 downto 0);
    output_voltage_cmd_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_voltage_unl_valid       : out std_logic;
    output_voltage_unl_ready       : in std_logic;
    output_voltage_unl_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0)
  );
end entity;

architecture Implementation of battery_status_output is
  -- signal voltage_inst_bcd_clk         : std_logic;
  signal voltage_inst_bcd_reset       : std_logic;

  -- signal voltage_inst_kcd_clk         : std_logic;
  signal voltage_inst_kcd_reset       : std_logic;

  signal voltage_inst_cmd_valid       : std_logic;
  signal voltage_inst_cmd_ready       : std_logic;
  signal voltage_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal voltage_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal voltage_inst_cmd_ctrl        : std_logic_vector(OUTPUT_VOLTAGE_BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal voltage_inst_cmd_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal voltage_inst_unl_valid       : std_logic;
  signal voltage_inst_unl_ready       : std_logic;
  signal voltage_inst_unl_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal voltage_inst_bus_wreq_valid  : std_logic;
  signal voltage_inst_bus_wreq_ready  : std_logic;
  signal voltage_inst_bus_wreq_addr   : std_logic_vector(OUTPUT_VOLTAGE_BUS_ADDR_WIDTH - 1 downto 0);
  signal voltage_inst_bus_wreq_len    : std_logic_vector(OUTPUT_VOLTAGE_BUS_LEN_WIDTH - 1 downto 0);
  signal voltage_inst_bus_wdat_valid  : std_logic;
  signal voltage_inst_bus_wdat_ready  : std_logic;
  signal voltage_inst_bus_wdat_data   : std_logic_vector(OUTPUT_VOLTAGE_BUS_DATA_WIDTH - 1 downto 0);
  signal voltage_inst_bus_wdat_strobe : std_logic_vector(OUTPUT_VOLTAGE_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal voltage_inst_bus_wdat_last   : std_logic;

  signal voltage_inst_in_valid        : std_logic_vector(1 downto 0);
  signal voltage_inst_in_ready        : std_logic_vector(1 downto 0);
  signal voltage_inst_in_data         : std_logic_vector(97 downto 0);
  signal voltage_inst_in_dvalid       : std_logic_vector(1 downto 0);
  signal voltage_inst_in_last         : std_logic_vector(1 downto 0);

begin
  voltage_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => OUTPUT_VOLTAGE_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => OUTPUT_VOLTAGE_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => OUTPUT_VOLTAGE_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => OUTPUT_VOLTAGE_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => OUTPUT_VOLTAGE_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "listprim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => voltage_inst_bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => voltage_inst_kcd_reset,
    cmd_valid       => voltage_inst_cmd_valid,
    cmd_ready       => voltage_inst_cmd_ready,
    cmd_firstIdx    => voltage_inst_cmd_firstIdx,
    cmd_lastIdx     => voltage_inst_cmd_lastIdx,
    cmd_ctrl        => voltage_inst_cmd_ctrl,
    cmd_tag         => voltage_inst_cmd_tag,
    unl_valid       => voltage_inst_unl_valid,
    unl_ready       => voltage_inst_unl_ready,
    unl_tag         => voltage_inst_unl_tag,
    bus_wreq_valid  => voltage_inst_bus_wreq_valid,
    bus_wreq_ready  => voltage_inst_bus_wreq_ready,
    bus_wreq_addr   => voltage_inst_bus_wreq_addr,
    bus_wreq_len    => voltage_inst_bus_wreq_len,
    bus_wdat_valid  => voltage_inst_bus_wdat_valid,
    bus_wdat_ready  => voltage_inst_bus_wdat_ready,
    bus_wdat_data   => voltage_inst_bus_wdat_data,
    bus_wdat_strobe => voltage_inst_bus_wdat_strobe,
    bus_wdat_last   => voltage_inst_bus_wdat_last,
    in_valid        => voltage_inst_in_valid,
    in_ready        => voltage_inst_in_ready,
    in_data         => voltage_inst_in_data,
    in_dvalid       => voltage_inst_in_dvalid,
    in_last         => voltage_inst_in_last
  );

  output_voltage_bus_wreq_valid      <= voltage_inst_bus_wreq_valid;
  voltage_inst_bus_wreq_ready        <= output_voltage_bus_wreq_ready;
  output_voltage_bus_wreq_addr       <= voltage_inst_bus_wreq_addr;
  output_voltage_bus_wreq_len        <= voltage_inst_bus_wreq_len;
  output_voltage_bus_wdat_valid      <= voltage_inst_bus_wdat_valid;
  voltage_inst_bus_wdat_ready        <= output_voltage_bus_wdat_ready;
  output_voltage_bus_wdat_data       <= voltage_inst_bus_wdat_data;
  output_voltage_bus_wdat_strobe     <= voltage_inst_bus_wdat_strobe;
  output_voltage_bus_wdat_last       <= voltage_inst_bus_wdat_last;

  output_voltage_unl_valid           <= voltage_inst_unl_valid;
  voltage_inst_unl_ready             <= output_voltage_unl_ready;
  output_voltage_unl_tag             <= voltage_inst_unl_tag;

  -- voltage_inst_bcd_clk               <= bcd_clk;
  voltage_inst_bcd_reset             <= bcd_reset;

  -- voltage_inst_kcd_clk               <= kcd_clk;
  voltage_inst_kcd_reset             <= kcd_reset;

  voltage_inst_cmd_valid             <= output_voltage_cmd_valid;
  output_voltage_cmd_ready           <= voltage_inst_cmd_ready;
  voltage_inst_cmd_firstIdx          <= output_voltage_cmd_firstIdx;
  voltage_inst_cmd_lastIdx           <= output_voltage_cmd_lastIdx;
  voltage_inst_cmd_ctrl              <= output_voltage_cmd_ctrl;
  voltage_inst_cmd_tag               <= output_voltage_cmd_tag;

  voltage_inst_in_valid(0)           <= output_voltage_valid;
  voltage_inst_in_valid(1)           <= output_voltage_item_valid;
  output_voltage_ready               <= voltage_inst_in_ready(0);
  output_voltage_item_ready          <= voltage_inst_in_ready(1);
  voltage_inst_in_data(31 downto 0)  <= output_voltage_length;
  voltage_inst_in_data(32 downto 32) <= output_voltage_count;
  voltage_inst_in_data(96 downto 33) <= output_voltage_item;
  voltage_inst_in_data(97 downto 97) <= output_voltage_item_count;
  voltage_inst_in_dvalid(0)          <= output_voltage_dvalid;
  voltage_inst_in_dvalid(1)          <= output_voltage_item_dvalid;
  voltage_inst_in_last(0)            <= output_voltage_last;
  voltage_inst_in_last(1)            <= output_voltage_item_last;

end architecture;