-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity battery_status_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk            : in std_logic;
    bcd_reset          : in std_logic;
    kcd_clk            : in std_logic;
    kcd_reset          : in std_logic;
    mmio_awvalid       : in std_logic;
    mmio_awready       : out std_logic;
    mmio_awaddr        : in std_logic_vector(31 downto 0);
    mmio_wvalid        : in std_logic;
    mmio_wready        : out std_logic;
    mmio_wdata         : in std_logic_vector(63 downto 0);
    mmio_wstrb         : in std_logic_vector(7 downto 0);
    mmio_bvalid        : out std_logic;
    mmio_bready        : in std_logic;
    mmio_bresp         : out std_logic_vector(1 downto 0);
    mmio_arvalid       : in std_logic;
    mmio_arready       : out std_logic;
    mmio_araddr        : in std_logic_vector(31 downto 0);
    mmio_rvalid        : out std_logic;
    mmio_rready        : in std_logic;
    mmio_rdata         : out std_logic_vector(63 downto 0);
    mmio_rresp         : out std_logic_vector(1 downto 0);
    rd_mst_rreq_valid  : out std_logic;
    rd_mst_rreq_ready  : in std_logic;
    rd_mst_rreq_addr   : out std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
    rd_mst_rreq_len    : out std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
    rd_mst_rdat_valid  : in std_logic;
    rd_mst_rdat_ready  : out std_logic;
    rd_mst_rdat_data   : in std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
    rd_mst_rdat_last   : in std_logic;
    wr_mst_wreq_valid  : out std_logic;
    wr_mst_wreq_ready  : in std_logic;
    wr_mst_wreq_addr   : out std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
    wr_mst_wreq_len    : out std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
    wr_mst_wdat_valid  : out std_logic;
    wr_mst_wdat_ready  : in std_logic;
    wr_mst_wdat_data   : out std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
    wr_mst_wdat_strobe : out std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
    wr_mst_wdat_last   : out std_logic;
    -- Platform completion handshake
    -- Assert req to indicate that the kernel is done, then ack will be strobed
    -- to indicate that the platform has finished propagating and publishing
    -- the write data.
    plat_complete_req  : out std_logic;
    plat_complete_ack  : in std_logic
  );
end entity;

architecture Implementation of battery_status_Mantle is
  component battery_status_Nucleus is
    generic (
      INDEX_WIDTH                   : integer := 32;
      TAG_WIDTH                     : integer := 1;
      INPUT_INPUT_BUS_ADDR_WIDTH    : integer := 64;
      OUTPUT_VOLTAGE_BUS_ADDR_WIDTH : integer := 64
    );
    port (
      kcd_clk                     : in std_logic;
      kcd_reset                   : in std_logic;
      mmio_awvalid                : in std_logic;
      mmio_awready                : out std_logic;
      mmio_awaddr                 : in std_logic_vector(31 downto 0);
      mmio_wvalid                 : in std_logic;
      mmio_wready                 : out std_logic;
      mmio_wdata                  : in std_logic_vector(63 downto 0);
      mmio_wstrb                  : in std_logic_vector(7 downto 0);
      mmio_bvalid                 : out std_logic;
      mmio_bready                 : in std_logic;
      mmio_bresp                  : out std_logic_vector(1 downto 0);
      mmio_arvalid                : in std_logic;
      mmio_arready                : out std_logic;
      mmio_araddr                 : in std_logic_vector(31 downto 0);
      mmio_rvalid                 : out std_logic;
      mmio_rready                 : in std_logic;
      mmio_rdata                  : out std_logic_vector(63 downto 0);
      mmio_rresp                  : out std_logic_vector(1 downto 0);
      input_input_valid           : in std_logic;
      input_input_ready           : out std_logic;
      input_input_dvalid          : in std_logic;
      input_input_last            : in std_logic;
      input_input                 : in std_logic_vector(63 downto 0);
      input_input_count           : in std_logic_vector(3 downto 0);
      input_input_unl_valid       : in std_logic;
      input_input_unl_ready       : out std_logic;
      input_input_unl_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      input_input_cmd_valid       : out std_logic;
      input_input_cmd_ready       : in std_logic;
      input_input_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      input_input_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      input_input_cmd_ctrl        : out std_logic_vector(INPUT_INPUT_BUS_ADDR_WIDTH - 1 downto 0);
      input_input_cmd_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      output_voltage_valid        : out std_logic;
      output_voltage_ready        : in std_logic;
      output_voltage_dvalid       : out std_logic;
      output_voltage_last         : out std_logic;
      output_voltage_length       : out std_logic_vector(31 downto 0);
      output_voltage_count        : out std_logic_vector(0 downto 0);
      output_voltage_item_valid   : out std_logic;
      output_voltage_item_ready   : in std_logic;
      output_voltage_item_dvalid  : out std_logic;
      output_voltage_item_last    : out std_logic;
      output_voltage_item         : out std_logic_vector(63 downto 0);
      output_voltage_item_count   : out std_logic_vector(0 downto 0);
      output_voltage_unl_valid    : in std_logic;
      output_voltage_unl_ready    : out std_logic;
      output_voltage_unl_tag      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      output_voltage_cmd_valid    : out std_logic;
      output_voltage_cmd_ready    : in std_logic;
      output_voltage_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      output_voltage_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      output_voltage_cmd_ctrl     : out std_logic_vector(OUTPUT_VOLTAGE_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      output_voltage_cmd_tag      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      plat_complete_req           : out std_logic;
      plat_complete_ack           : in std_logic
    );
  end component;

  component battery_status_input is
    generic (
      INDEX_WIDTH                    : integer := 32;
      TAG_WIDTH                      : integer := 1;
      INPUT_INPUT_BUS_ADDR_WIDTH     : integer := 64;
      INPUT_INPUT_BUS_DATA_WIDTH     : integer := 512;
      INPUT_INPUT_BUS_LEN_WIDTH      : integer := 8;
      INPUT_INPUT_BUS_BURST_STEP_LEN : integer := 1;
      INPUT_INPUT_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                    : in std_logic;
      bcd_reset                  : in std_logic;
      kcd_clk                    : in std_logic;
      kcd_reset                  : in std_logic;
      input_input_valid          : out std_logic;
      input_input_ready          : in std_logic;
      input_input_dvalid         : out std_logic;
      input_input_last           : out std_logic;
      input_input                : out std_logic_vector(63 downto 0);
      input_input_count          : out std_logic_vector(3 downto 0);
      input_input_bus_rreq_valid : out std_logic;
      input_input_bus_rreq_ready : in std_logic;
      input_input_bus_rreq_addr  : out std_logic_vector(INPUT_INPUT_BUS_ADDR_WIDTH - 1 downto 0);
      input_input_bus_rreq_len   : out std_logic_vector(INPUT_INPUT_BUS_LEN_WIDTH - 1 downto 0);
      input_input_bus_rdat_valid : in std_logic;
      input_input_bus_rdat_ready : out std_logic;
      input_input_bus_rdat_data  : in std_logic_vector(INPUT_INPUT_BUS_DATA_WIDTH - 1 downto 0);
      input_input_bus_rdat_last  : in std_logic;
      input_input_cmd_valid      : in std_logic;
      input_input_cmd_ready      : out std_logic;
      input_input_cmd_firstIdx   : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      input_input_cmd_lastIdx    : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      input_input_cmd_ctrl       : in std_logic_vector(INPUT_INPUT_BUS_ADDR_WIDTH - 1 downto 0);
      input_input_cmd_tag        : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      input_input_unl_valid      : out std_logic;
      input_input_unl_ready      : in std_logic;
      input_input_unl_tag        : out std_logic_vector(TAG_WIDTH - 1 downto 0)
    );
  end component;

  component battery_status_output is
    generic (
      INDEX_WIDTH                       : integer := 32;
      TAG_WIDTH                         : integer := 1;
      OUTPUT_VOLTAGE_BUS_ADDR_WIDTH     : integer := 64;
      OUTPUT_VOLTAGE_BUS_DATA_WIDTH     : integer := 512;
      OUTPUT_VOLTAGE_BUS_LEN_WIDTH      : integer := 8;
      OUTPUT_VOLTAGE_BUS_BURST_STEP_LEN : integer := 1;
      OUTPUT_VOLTAGE_BUS_BURST_MAX_LEN  : integer := 16
    );
    port (
      bcd_clk                        : in std_logic;
      bcd_reset                      : in std_logic;
      kcd_clk                        : in std_logic;
      kcd_reset                      : in std_logic;
      output_voltage_valid           : in std_logic;
      output_voltage_ready           : out std_logic;
      output_voltage_dvalid          : in std_logic;
      output_voltage_last            : in std_logic;
      output_voltage_length          : in std_logic_vector(31 downto 0);
      output_voltage_count           : in std_logic_vector(0 downto 0);
      output_voltage_item_valid      : in std_logic;
      output_voltage_item_ready      : out std_logic;
      output_voltage_item_dvalid     : in std_logic;
      output_voltage_item_last       : in std_logic;
      output_voltage_item            : in std_logic_vector(63 downto 0);
      output_voltage_item_count      : in std_logic_vector(0 downto 0);
      output_voltage_bus_wreq_valid  : out std_logic;
      output_voltage_bus_wreq_ready  : in std_logic;
      output_voltage_bus_wreq_addr   : out std_logic_vector(OUTPUT_VOLTAGE_BUS_ADDR_WIDTH - 1 downto 0);
      output_voltage_bus_wreq_len    : out std_logic_vector(OUTPUT_VOLTAGE_BUS_LEN_WIDTH - 1 downto 0);
      output_voltage_bus_wdat_valid  : out std_logic;
      output_voltage_bus_wdat_ready  : in std_logic;
      output_voltage_bus_wdat_data   : out std_logic_vector(OUTPUT_VOLTAGE_BUS_DATA_WIDTH - 1 downto 0);
      output_voltage_bus_wdat_strobe : out std_logic_vector(OUTPUT_VOLTAGE_BUS_DATA_WIDTH/8 - 1 downto 0);
      output_voltage_bus_wdat_last   : out std_logic;
      output_voltage_cmd_valid       : in std_logic;
      output_voltage_cmd_ready       : out std_logic;
      output_voltage_cmd_firstIdx    : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      output_voltage_cmd_lastIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      output_voltage_cmd_ctrl        : in std_logic_vector(OUTPUT_VOLTAGE_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      output_voltage_cmd_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      output_voltage_unl_valid       : out std_logic;
      output_voltage_unl_ready       : in std_logic;
      output_voltage_unl_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0)
    );
  end component;

  signal battery_status_Nucleus_inst_kcd_clk                       : std_logic;
  signal battery_status_Nucleus_inst_kcd_reset                     : std_logic;

  signal battery_status_Nucleus_inst_mmio_awvalid                  : std_logic;
  signal battery_status_Nucleus_inst_mmio_awready                  : std_logic;
  signal battery_status_Nucleus_inst_mmio_awaddr                   : std_logic_vector(31 downto 0);
  signal battery_status_Nucleus_inst_mmio_wvalid                   : std_logic;
  signal battery_status_Nucleus_inst_mmio_wready                   : std_logic;
  signal battery_status_Nucleus_inst_mmio_wdata                    : std_logic_vector(63 downto 0);
  signal battery_status_Nucleus_inst_mmio_wstrb                    : std_logic_vector(7 downto 0);
  signal battery_status_Nucleus_inst_mmio_bvalid                   : std_logic;
  signal battery_status_Nucleus_inst_mmio_bready                   : std_logic;
  signal battery_status_Nucleus_inst_mmio_bresp                    : std_logic_vector(1 downto 0);
  signal battery_status_Nucleus_inst_mmio_arvalid                  : std_logic;
  signal battery_status_Nucleus_inst_mmio_arready                  : std_logic;
  signal battery_status_Nucleus_inst_mmio_araddr                   : std_logic_vector(31 downto 0);
  signal battery_status_Nucleus_inst_mmio_rvalid                   : std_logic;
  signal battery_status_Nucleus_inst_mmio_rready                   : std_logic;
  signal battery_status_Nucleus_inst_mmio_rdata                    : std_logic_vector(63 downto 0);
  signal battery_status_Nucleus_inst_mmio_rresp                    : std_logic_vector(1 downto 0);

  signal battery_status_Nucleus_inst_input_input_valid             : std_logic;
  signal battery_status_Nucleus_inst_input_input_ready             : std_logic;
  signal battery_status_Nucleus_inst_input_input_dvalid            : std_logic;
  signal battery_status_Nucleus_inst_input_input_last              : std_logic;
  signal battery_status_Nucleus_inst_input_input                   : std_logic_vector(63 downto 0);
  signal battery_status_Nucleus_inst_input_input_count             : std_logic_vector(3 downto 0);

  signal battery_status_Nucleus_inst_input_input_unl_valid         : std_logic;
  signal battery_status_Nucleus_inst_input_input_unl_ready         : std_logic;
  signal battery_status_Nucleus_inst_input_input_unl_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal battery_status_Nucleus_inst_input_input_cmd_valid         : std_logic;
  signal battery_status_Nucleus_inst_input_input_cmd_ready         : std_logic;
  signal battery_status_Nucleus_inst_input_input_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_Nucleus_inst_input_input_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_Nucleus_inst_input_input_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal battery_status_Nucleus_inst_input_input_cmd_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal battery_status_Nucleus_inst_output_voltage_valid          : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_ready          : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_dvalid         : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_last           : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_length         : std_logic_vector(31 downto 0);
  signal battery_status_Nucleus_inst_output_voltage_count          : std_logic_vector(0 downto 0);
  signal battery_status_Nucleus_inst_output_voltage_item_valid     : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_item_ready     : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_item_dvalid    : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_item_last      : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_item           : std_logic_vector(63 downto 0);
  signal battery_status_Nucleus_inst_output_voltage_item_count     : std_logic_vector(0 downto 0);

  signal battery_status_Nucleus_inst_output_voltage_unl_valid      : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_unl_ready      : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_unl_tag        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal battery_status_Nucleus_inst_output_voltage_cmd_valid      : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_cmd_ready      : std_logic;
  signal battery_status_Nucleus_inst_output_voltage_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_Nucleus_inst_output_voltage_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_Nucleus_inst_output_voltage_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal battery_status_Nucleus_inst_output_voltage_cmd_tag        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal battery_status_input_inst_bcd_clk                         : std_logic;
  signal battery_status_input_inst_bcd_reset                       : std_logic;

  signal battery_status_input_inst_kcd_clk                         : std_logic;
  signal battery_status_input_inst_kcd_reset                       : std_logic;

  signal battery_status_input_inst_input_input_valid               : std_logic;
  signal battery_status_input_inst_input_input_ready               : std_logic;
  signal battery_status_input_inst_input_input_dvalid              : std_logic;
  signal battery_status_input_inst_input_input_last                : std_logic;
  signal battery_status_input_inst_input_input                     : std_logic_vector(63 downto 0);
  signal battery_status_input_inst_input_input_count               : std_logic_vector(3 downto 0);

  signal battery_status_input_inst_input_input_bus_rreq_valid      : std_logic;
  signal battery_status_input_inst_input_input_bus_rreq_ready      : std_logic;
  signal battery_status_input_inst_input_input_bus_rreq_addr       : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal battery_status_input_inst_input_input_bus_rreq_len        : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal battery_status_input_inst_input_input_bus_rdat_valid      : std_logic;
  signal battery_status_input_inst_input_input_bus_rdat_ready      : std_logic;
  signal battery_status_input_inst_input_input_bus_rdat_data       : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal battery_status_input_inst_input_input_bus_rdat_last       : std_logic;

  signal battery_status_input_inst_input_input_cmd_valid           : std_logic;
  signal battery_status_input_inst_input_input_cmd_ready           : std_logic;
  signal battery_status_input_inst_input_input_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_input_inst_input_input_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_input_inst_input_input_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal battery_status_input_inst_input_input_cmd_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal battery_status_input_inst_input_input_unl_valid           : std_logic;
  signal battery_status_input_inst_input_input_unl_ready           : std_logic;
  signal battery_status_input_inst_input_input_unl_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal battery_status_output_inst_bcd_clk                        : std_logic;
  signal battery_status_output_inst_bcd_reset                      : std_logic;

  signal battery_status_output_inst_kcd_clk                        : std_logic;
  signal battery_status_output_inst_kcd_reset                      : std_logic;

  signal battery_status_output_inst_output_voltage_valid           : std_logic;
  signal battery_status_output_inst_output_voltage_ready           : std_logic;
  signal battery_status_output_inst_output_voltage_dvalid          : std_logic;
  signal battery_status_output_inst_output_voltage_last            : std_logic;
  signal battery_status_output_inst_output_voltage_length          : std_logic_vector(31 downto 0);
  signal battery_status_output_inst_output_voltage_count           : std_logic_vector(0 downto 0);
  signal battery_status_output_inst_output_voltage_item_valid      : std_logic;
  signal battery_status_output_inst_output_voltage_item_ready      : std_logic;
  signal battery_status_output_inst_output_voltage_item_dvalid     : std_logic;
  signal battery_status_output_inst_output_voltage_item_last       : std_logic;
  signal battery_status_output_inst_output_voltage_item            : std_logic_vector(63 downto 0);
  signal battery_status_output_inst_output_voltage_item_count      : std_logic_vector(0 downto 0);

  signal battery_status_output_inst_output_voltage_bus_wreq_valid  : std_logic;
  signal battery_status_output_inst_output_voltage_bus_wreq_ready  : std_logic;
  signal battery_status_output_inst_output_voltage_bus_wreq_addr   : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal battery_status_output_inst_output_voltage_bus_wreq_len    : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal battery_status_output_inst_output_voltage_bus_wdat_valid  : std_logic;
  signal battery_status_output_inst_output_voltage_bus_wdat_ready  : std_logic;
  signal battery_status_output_inst_output_voltage_bus_wdat_data   : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal battery_status_output_inst_output_voltage_bus_wdat_strobe : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal battery_status_output_inst_output_voltage_bus_wdat_last   : std_logic;

  signal battery_status_output_inst_output_voltage_cmd_valid       : std_logic;
  signal battery_status_output_inst_output_voltage_cmd_ready       : std_logic;
  signal battery_status_output_inst_output_voltage_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_output_inst_output_voltage_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal battery_status_output_inst_output_voltage_cmd_ctrl        : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal battery_status_output_inst_output_voltage_cmd_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal battery_status_output_inst_output_voltage_unl_valid       : std_logic;
  signal battery_status_output_inst_output_voltage_unl_ready       : std_logic;
  signal battery_status_output_inst_output_voltage_unl_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal RDAW64DW512LW8BS1BM16_inst_bcd_clk                        : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_bcd_reset                      : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_len                   : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready                 : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_data                  : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_last                  : std_logic;

  signal WRAW64DW512LW8BS1BM16_inst_bcd_clk                        : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_bcd_reset                      : std_logic;

  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_len                   : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready                 : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_data                  : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe                : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_last                  : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid                 : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready                 : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len                   : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid                 : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready                 : std_logic_vector(0 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data                  : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last                  : std_logic_vector(0 downto 0);

  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid                 : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready                 : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len                   : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid                 : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready                 : std_logic_vector(0 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data                  : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe                : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last                  : std_logic_vector(0 downto 0);

begin
  battery_status_Nucleus_inst : battery_status_Nucleus
  generic map(
    INDEX_WIDTH                   => INDEX_WIDTH,
    TAG_WIDTH                     => TAG_WIDTH,
    INPUT_INPUT_BUS_ADDR_WIDTH    => BUS_ADDR_WIDTH,
    OUTPUT_VOLTAGE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH
  )
  port map(
    kcd_clk                     => battery_status_Nucleus_inst_kcd_clk,
    kcd_reset                   => battery_status_Nucleus_inst_kcd_reset,
    mmio_awvalid                => battery_status_Nucleus_inst_mmio_awvalid,
    mmio_awready                => battery_status_Nucleus_inst_mmio_awready,
    mmio_awaddr                 => battery_status_Nucleus_inst_mmio_awaddr,
    mmio_wvalid                 => battery_status_Nucleus_inst_mmio_wvalid,
    mmio_wready                 => battery_status_Nucleus_inst_mmio_wready,
    mmio_wdata                  => battery_status_Nucleus_inst_mmio_wdata,
    mmio_wstrb                  => battery_status_Nucleus_inst_mmio_wstrb,
    mmio_bvalid                 => battery_status_Nucleus_inst_mmio_bvalid,
    mmio_bready                 => battery_status_Nucleus_inst_mmio_bready,
    mmio_bresp                  => battery_status_Nucleus_inst_mmio_bresp,
    mmio_arvalid                => battery_status_Nucleus_inst_mmio_arvalid,
    mmio_arready                => battery_status_Nucleus_inst_mmio_arready,
    mmio_araddr                 => battery_status_Nucleus_inst_mmio_araddr,
    mmio_rvalid                 => battery_status_Nucleus_inst_mmio_rvalid,
    mmio_rready                 => battery_status_Nucleus_inst_mmio_rready,
    mmio_rdata                  => battery_status_Nucleus_inst_mmio_rdata,
    mmio_rresp                  => battery_status_Nucleus_inst_mmio_rresp,
    input_input_valid           => battery_status_Nucleus_inst_input_input_valid,
    input_input_ready           => battery_status_Nucleus_inst_input_input_ready,
    input_input_dvalid          => battery_status_Nucleus_inst_input_input_dvalid,
    input_input_last            => battery_status_Nucleus_inst_input_input_last,
    input_input                 => battery_status_Nucleus_inst_input_input,
    input_input_count           => battery_status_Nucleus_inst_input_input_count,
    input_input_unl_valid       => battery_status_Nucleus_inst_input_input_unl_valid,
    input_input_unl_ready       => battery_status_Nucleus_inst_input_input_unl_ready,
    input_input_unl_tag         => battery_status_Nucleus_inst_input_input_unl_tag,
    input_input_cmd_valid       => battery_status_Nucleus_inst_input_input_cmd_valid,
    input_input_cmd_ready       => battery_status_Nucleus_inst_input_input_cmd_ready,
    input_input_cmd_firstIdx    => battery_status_Nucleus_inst_input_input_cmd_firstIdx,
    input_input_cmd_lastIdx     => battery_status_Nucleus_inst_input_input_cmd_lastIdx,
    input_input_cmd_ctrl        => battery_status_Nucleus_inst_input_input_cmd_ctrl,
    input_input_cmd_tag         => battery_status_Nucleus_inst_input_input_cmd_tag,
    output_voltage_valid        => battery_status_Nucleus_inst_output_voltage_valid,
    output_voltage_ready        => battery_status_Nucleus_inst_output_voltage_ready,
    output_voltage_dvalid       => battery_status_Nucleus_inst_output_voltage_dvalid,
    output_voltage_last         => battery_status_Nucleus_inst_output_voltage_last,
    output_voltage_length       => battery_status_Nucleus_inst_output_voltage_length,
    output_voltage_count        => battery_status_Nucleus_inst_output_voltage_count,
    output_voltage_item_valid   => battery_status_Nucleus_inst_output_voltage_item_valid,
    output_voltage_item_ready   => battery_status_Nucleus_inst_output_voltage_item_ready,
    output_voltage_item_dvalid  => battery_status_Nucleus_inst_output_voltage_item_dvalid,
    output_voltage_item_last    => battery_status_Nucleus_inst_output_voltage_item_last,
    output_voltage_item         => battery_status_Nucleus_inst_output_voltage_item,
    output_voltage_item_count   => battery_status_Nucleus_inst_output_voltage_item_count,
    output_voltage_unl_valid    => battery_status_Nucleus_inst_output_voltage_unl_valid,
    output_voltage_unl_ready    => battery_status_Nucleus_inst_output_voltage_unl_ready,
    output_voltage_unl_tag      => battery_status_Nucleus_inst_output_voltage_unl_tag,
    output_voltage_cmd_valid    => battery_status_Nucleus_inst_output_voltage_cmd_valid,
    output_voltage_cmd_ready    => battery_status_Nucleus_inst_output_voltage_cmd_ready,
    output_voltage_cmd_firstIdx => battery_status_Nucleus_inst_output_voltage_cmd_firstIdx,
    output_voltage_cmd_lastIdx  => battery_status_Nucleus_inst_output_voltage_cmd_lastIdx,
    output_voltage_cmd_ctrl     => battery_status_Nucleus_inst_output_voltage_cmd_ctrl,
    output_voltage_cmd_tag      => battery_status_Nucleus_inst_output_voltage_cmd_tag,
    plat_complete_ack           => plat_complete_ack,
    plat_complete_req           => plat_complete_req
  );

  battery_status_input_inst : battery_status_input
  generic map(
    INDEX_WIDTH                    => INDEX_WIDTH,
    TAG_WIDTH                      => TAG_WIDTH,
    INPUT_INPUT_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
    INPUT_INPUT_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
    INPUT_INPUT_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
    INPUT_INPUT_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    INPUT_INPUT_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
  )
  port map(
    bcd_clk                    => battery_status_input_inst_bcd_clk,
    bcd_reset                  => battery_status_input_inst_bcd_reset,
    kcd_clk                    => battery_status_input_inst_kcd_clk,
    kcd_reset                  => battery_status_input_inst_kcd_reset,
    input_input_valid          => battery_status_input_inst_input_input_valid,
    input_input_ready          => battery_status_input_inst_input_input_ready,
    input_input_dvalid         => battery_status_input_inst_input_input_dvalid,
    input_input_last           => battery_status_input_inst_input_input_last,
    input_input                => battery_status_input_inst_input_input,
    input_input_count          => battery_status_input_inst_input_input_count,
    input_input_bus_rreq_valid => battery_status_input_inst_input_input_bus_rreq_valid,
    input_input_bus_rreq_ready => battery_status_input_inst_input_input_bus_rreq_ready,
    input_input_bus_rreq_addr  => battery_status_input_inst_input_input_bus_rreq_addr,
    input_input_bus_rreq_len   => battery_status_input_inst_input_input_bus_rreq_len,
    input_input_bus_rdat_valid => battery_status_input_inst_input_input_bus_rdat_valid,
    input_input_bus_rdat_ready => battery_status_input_inst_input_input_bus_rdat_ready,
    input_input_bus_rdat_data  => battery_status_input_inst_input_input_bus_rdat_data,
    input_input_bus_rdat_last  => battery_status_input_inst_input_input_bus_rdat_last,
    input_input_cmd_valid      => battery_status_input_inst_input_input_cmd_valid,
    input_input_cmd_ready      => battery_status_input_inst_input_input_cmd_ready,
    input_input_cmd_firstIdx   => battery_status_input_inst_input_input_cmd_firstIdx,
    input_input_cmd_lastIdx    => battery_status_input_inst_input_input_cmd_lastIdx,
    input_input_cmd_ctrl       => battery_status_input_inst_input_input_cmd_ctrl,
    input_input_cmd_tag        => battery_status_input_inst_input_input_cmd_tag,
    input_input_unl_valid      => battery_status_input_inst_input_input_unl_valid,
    input_input_unl_ready      => battery_status_input_inst_input_input_unl_ready,
    input_input_unl_tag        => battery_status_input_inst_input_input_unl_tag
  );

  battery_status_output_inst : battery_status_output
  generic map(
    INDEX_WIDTH                       => INDEX_WIDTH,
    TAG_WIDTH                         => TAG_WIDTH,
    OUTPUT_VOLTAGE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
    OUTPUT_VOLTAGE_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
    OUTPUT_VOLTAGE_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
    OUTPUT_VOLTAGE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    OUTPUT_VOLTAGE_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN
  )
  port map(
    bcd_clk                        => battery_status_output_inst_bcd_clk,
    bcd_reset                      => battery_status_output_inst_bcd_reset,
    kcd_clk                        => battery_status_output_inst_kcd_clk,
    kcd_reset                      => battery_status_output_inst_kcd_reset,
    output_voltage_valid           => battery_status_output_inst_output_voltage_valid,
    output_voltage_ready           => battery_status_output_inst_output_voltage_ready,
    output_voltage_dvalid          => battery_status_output_inst_output_voltage_dvalid,
    output_voltage_last            => battery_status_output_inst_output_voltage_last,
    output_voltage_length          => battery_status_output_inst_output_voltage_length,
    output_voltage_count           => battery_status_output_inst_output_voltage_count,
    output_voltage_item_valid      => battery_status_output_inst_output_voltage_item_valid,
    output_voltage_item_ready      => battery_status_output_inst_output_voltage_item_ready,
    output_voltage_item_dvalid     => battery_status_output_inst_output_voltage_item_dvalid,
    output_voltage_item_last       => battery_status_output_inst_output_voltage_item_last,
    output_voltage_item            => battery_status_output_inst_output_voltage_item,
    output_voltage_item_count      => battery_status_output_inst_output_voltage_item_count,
    output_voltage_bus_wreq_valid  => battery_status_output_inst_output_voltage_bus_wreq_valid,
    output_voltage_bus_wreq_ready  => battery_status_output_inst_output_voltage_bus_wreq_ready,
    output_voltage_bus_wreq_addr   => battery_status_output_inst_output_voltage_bus_wreq_addr,
    output_voltage_bus_wreq_len    => battery_status_output_inst_output_voltage_bus_wreq_len,
    output_voltage_bus_wdat_valid  => battery_status_output_inst_output_voltage_bus_wdat_valid,
    output_voltage_bus_wdat_ready  => battery_status_output_inst_output_voltage_bus_wdat_ready,
    output_voltage_bus_wdat_data   => battery_status_output_inst_output_voltage_bus_wdat_data,
    output_voltage_bus_wdat_strobe => battery_status_output_inst_output_voltage_bus_wdat_strobe,
    output_voltage_bus_wdat_last   => battery_status_output_inst_output_voltage_bus_wdat_last,
    output_voltage_cmd_valid       => battery_status_output_inst_output_voltage_cmd_valid,
    output_voltage_cmd_ready       => battery_status_output_inst_output_voltage_cmd_ready,
    output_voltage_cmd_firstIdx    => battery_status_output_inst_output_voltage_cmd_firstIdx,
    output_voltage_cmd_lastIdx     => battery_status_output_inst_output_voltage_cmd_lastIdx,
    output_voltage_cmd_ctrl        => battery_status_output_inst_output_voltage_cmd_ctrl,
    output_voltage_cmd_tag         => battery_status_output_inst_output_voltage_cmd_tag,
    output_voltage_unl_valid       => battery_status_output_inst_output_voltage_unl_valid,
    output_voltage_unl_ready       => battery_status_output_inst_output_voltage_unl_ready,
    output_voltage_unl_tag         => battery_status_output_inst_output_voltage_unl_tag
  );

  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
  generic map(
    BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
    BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
    NUM_SLAVE_PORTS => 1,
    ARB_METHOD      => "RR-STICKY",
    MAX_OUTSTANDING => 4,
    RAM_CONFIG      => "",
    SLV_REQ_SLICES  => true,
    MST_REQ_SLICE   => true,
    MST_DAT_SLICE   => true,
    SLV_DAT_SLICES  => true
  )
  port map(
    bcd_clk        => RDAW64DW512LW8BS1BM16_inst_bcd_clk,
    bcd_reset      => RDAW64DW512LW8BS1BM16_inst_bcd_reset,
    mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
    mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
    mst_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
    mst_rreq_len   => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
    mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
    mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
    mst_rdat_data  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
    mst_rdat_last  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
    bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
    bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
    bsv_rreq_len   => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
    bsv_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
    bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
    bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
    bsv_rdat_last  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
    bsv_rdat_data  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
  );

  WRAW64DW512LW8BS1BM16_inst : BusWriteArbiterVec
  generic map(
    BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
    BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
    NUM_SLAVE_PORTS => 1,
    ARB_METHOD      => "RR-STICKY",
    MAX_OUTSTANDING => 4,
    RAM_CONFIG      => "",
    SLV_REQ_SLICES  => true,
    MST_REQ_SLICE   => true,
    MST_DAT_SLICE   => true,
    SLV_DAT_SLICES  => true
  )
  port map(
    bcd_clk         => WRAW64DW512LW8BS1BM16_inst_bcd_clk,
    bcd_reset       => WRAW64DW512LW8BS1BM16_inst_bcd_reset,
    mst_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid,
    mst_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready,
    mst_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr,
    mst_wreq_len    => WRAW64DW512LW8BS1BM16_inst_mst_wreq_len,
    mst_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid,
    mst_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready,
    mst_wdat_data   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_data,
    mst_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe,
    mst_wdat_last   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_last,
    bsv_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid,
    bsv_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready,
    bsv_wreq_len    => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len,
    bsv_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr,
    bsv_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid,
    bsv_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe,
    bsv_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready,
    bsv_wdat_last   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last,
    bsv_wdat_data   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data
  );

  rd_mst_rreq_valid                                                         <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready                                 <= rd_mst_rreq_ready;
  rd_mst_rreq_addr                                                          <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len                                                           <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid                                 <= rd_mst_rdat_valid;
  rd_mst_rdat_ready                                                         <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data                                  <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last                                  <= rd_mst_rdat_last;

  wr_mst_wreq_valid                                                         <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready                                 <= wr_mst_wreq_ready;
  wr_mst_wreq_addr                                                          <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr;
  wr_mst_wreq_len                                                           <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_len;
  wr_mst_wdat_valid                                                         <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready                                 <= wr_mst_wdat_ready;
  wr_mst_wdat_data                                                          <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_data;
  wr_mst_wdat_strobe                                                        <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe;
  wr_mst_wdat_last                                                          <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_last;

  battery_status_Nucleus_inst_kcd_clk                                       <= kcd_clk;
  battery_status_Nucleus_inst_kcd_reset                                     <= kcd_reset;

  battery_status_Nucleus_inst_mmio_awvalid                                  <= mmio_awvalid;
  mmio_awready                                                              <= battery_status_Nucleus_inst_mmio_awready;
  battery_status_Nucleus_inst_mmio_awaddr                                   <= mmio_awaddr;
  battery_status_Nucleus_inst_mmio_wvalid                                   <= mmio_wvalid;
  mmio_wready                                                               <= battery_status_Nucleus_inst_mmio_wready;
  battery_status_Nucleus_inst_mmio_wdata                                    <= mmio_wdata;
  battery_status_Nucleus_inst_mmio_wstrb                                    <= mmio_wstrb;
  mmio_bvalid                                                               <= battery_status_Nucleus_inst_mmio_bvalid;
  battery_status_Nucleus_inst_mmio_bready                                   <= mmio_bready;
  mmio_bresp                                                                <= battery_status_Nucleus_inst_mmio_bresp;
  battery_status_Nucleus_inst_mmio_arvalid                                  <= mmio_arvalid;
  mmio_arready                                                              <= battery_status_Nucleus_inst_mmio_arready;
  battery_status_Nucleus_inst_mmio_araddr                                   <= mmio_araddr;
  mmio_rvalid                                                               <= battery_status_Nucleus_inst_mmio_rvalid;
  battery_status_Nucleus_inst_mmio_rready                                   <= mmio_rready;
  mmio_rdata                                                                <= battery_status_Nucleus_inst_mmio_rdata;
  mmio_rresp                                                                <= battery_status_Nucleus_inst_mmio_rresp;

  battery_status_Nucleus_inst_input_input_valid                             <= battery_status_input_inst_input_input_valid;
  battery_status_input_inst_input_input_ready                               <= battery_status_Nucleus_inst_input_input_ready;
  battery_status_Nucleus_inst_input_input_dvalid                            <= battery_status_input_inst_input_input_dvalid;
  battery_status_Nucleus_inst_input_input_last                              <= battery_status_input_inst_input_input_last;
  battery_status_Nucleus_inst_input_input                                   <= battery_status_input_inst_input_input;
  battery_status_Nucleus_inst_input_input_count                             <= battery_status_input_inst_input_input_count;

  battery_status_Nucleus_inst_input_input_unl_valid                         <= battery_status_input_inst_input_input_unl_valid;
  battery_status_input_inst_input_input_unl_ready                           <= battery_status_Nucleus_inst_input_input_unl_ready;
  battery_status_Nucleus_inst_input_input_unl_tag                           <= battery_status_input_inst_input_input_unl_tag;

  battery_status_Nucleus_inst_output_voltage_unl_valid                      <= battery_status_output_inst_output_voltage_unl_valid;
  battery_status_output_inst_output_voltage_unl_ready                       <= battery_status_Nucleus_inst_output_voltage_unl_ready;
  battery_status_Nucleus_inst_output_voltage_unl_tag                        <= battery_status_output_inst_output_voltage_unl_tag;

  battery_status_input_inst_bcd_clk                                         <= bcd_clk;
  battery_status_input_inst_bcd_reset                                       <= bcd_reset;

  battery_status_input_inst_kcd_clk                                         <= kcd_clk;
  battery_status_input_inst_kcd_reset                                       <= kcd_reset;

  battery_status_input_inst_input_input_cmd_valid                           <= battery_status_Nucleus_inst_input_input_cmd_valid;
  battery_status_Nucleus_inst_input_input_cmd_ready                         <= battery_status_input_inst_input_input_cmd_ready;
  battery_status_input_inst_input_input_cmd_firstIdx                        <= battery_status_Nucleus_inst_input_input_cmd_firstIdx;
  battery_status_input_inst_input_input_cmd_lastIdx                         <= battery_status_Nucleus_inst_input_input_cmd_lastIdx;
  battery_status_input_inst_input_input_cmd_ctrl                            <= battery_status_Nucleus_inst_input_input_cmd_ctrl;
  battery_status_input_inst_input_input_cmd_tag                             <= battery_status_Nucleus_inst_input_input_cmd_tag;

  battery_status_output_inst_bcd_clk                                        <= bcd_clk;
  battery_status_output_inst_bcd_reset                                      <= bcd_reset;

  battery_status_output_inst_kcd_clk                                        <= kcd_clk;
  battery_status_output_inst_kcd_reset                                      <= kcd_reset;

  battery_status_output_inst_output_voltage_valid                           <= battery_status_Nucleus_inst_output_voltage_valid;
  battery_status_Nucleus_inst_output_voltage_ready                          <= battery_status_output_inst_output_voltage_ready;
  battery_status_output_inst_output_voltage_dvalid                          <= battery_status_Nucleus_inst_output_voltage_dvalid;
  battery_status_output_inst_output_voltage_last                            <= battery_status_Nucleus_inst_output_voltage_last;
  battery_status_output_inst_output_voltage_length                          <= battery_status_Nucleus_inst_output_voltage_length;
  battery_status_output_inst_output_voltage_count                           <= battery_status_Nucleus_inst_output_voltage_count;
  battery_status_output_inst_output_voltage_item_valid                      <= battery_status_Nucleus_inst_output_voltage_item_valid;
  battery_status_Nucleus_inst_output_voltage_item_ready                     <= battery_status_output_inst_output_voltage_item_ready;
  battery_status_output_inst_output_voltage_item_dvalid                     <= battery_status_Nucleus_inst_output_voltage_item_dvalid;
  battery_status_output_inst_output_voltage_item_last                       <= battery_status_Nucleus_inst_output_voltage_item_last;
  battery_status_output_inst_output_voltage_item                            <= battery_status_Nucleus_inst_output_voltage_item;
  battery_status_output_inst_output_voltage_item_count                      <= battery_status_Nucleus_inst_output_voltage_item_count;

  battery_status_output_inst_output_voltage_cmd_valid                       <= battery_status_Nucleus_inst_output_voltage_cmd_valid;
  battery_status_Nucleus_inst_output_voltage_cmd_ready                      <= battery_status_output_inst_output_voltage_cmd_ready;
  battery_status_output_inst_output_voltage_cmd_firstIdx                    <= battery_status_Nucleus_inst_output_voltage_cmd_firstIdx;
  battery_status_output_inst_output_voltage_cmd_lastIdx                     <= battery_status_Nucleus_inst_output_voltage_cmd_lastIdx;
  battery_status_output_inst_output_voltage_cmd_ctrl                        <= battery_status_Nucleus_inst_output_voltage_cmd_ctrl;
  battery_status_output_inst_output_voltage_cmd_tag                         <= battery_status_Nucleus_inst_output_voltage_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bcd_clk                                        <= bcd_clk;
  RDAW64DW512LW8BS1BM16_inst_bcd_reset                                      <= bcd_reset;

  WRAW64DW512LW8BS1BM16_inst_bcd_clk                                        <= bcd_clk;
  WRAW64DW512LW8BS1BM16_inst_bcd_reset                                      <= bcd_reset;

  battery_status_input_inst_input_input_bus_rreq_ready                      <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  battery_status_input_inst_input_input_bus_rdat_valid                      <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  battery_status_input_inst_input_input_bus_rdat_last                       <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  battery_status_input_inst_input_input_bus_rdat_data                       <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH - 1 downto 0);
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0)                              <= battery_status_input_inst_input_input_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH - 1 downto 0)       <= battery_status_input_inst_input_input_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH - 1 downto 0)     <= battery_status_input_inst_input_input_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0)                              <= battery_status_input_inst_input_input_bus_rdat_ready;

  battery_status_output_inst_output_voltage_bus_wreq_ready                  <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(0);
  battery_status_output_inst_output_voltage_bus_wdat_ready                  <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(0);
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(0)                              <= battery_status_output_inst_output_voltage_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH - 1 downto 0)       <= battery_status_output_inst_output_voltage_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH - 1 downto 0)     <= battery_status_output_inst_output_voltage_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(0)                              <= battery_status_output_inst_output_voltage_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 - 1 downto 0) <= battery_status_output_inst_output_voltage_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(0)                               <= battery_status_output_inst_output_voltage_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH - 1 downto 0)     <= battery_status_output_inst_output_voltage_bus_wdat_data;

end architecture;