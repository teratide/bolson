-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.battery_status_pkg.all;
use work.Stream_pkg.all;

entity battery_status_2 is
  generic (
    INDEX_WIDTH : integer := 32;
    TAG_WIDTH   : integer := 1
  );
  port (
    kcd_clk                       : in std_logic;
    kcd_reset                     : in std_logic;
    input_1_input_valid           : in std_logic;
    input_1_input_ready           : out std_logic;
    input_1_input_dvalid          : in std_logic;
    input_1_input_last            : in std_logic;
    input_1_input                 : in std_logic_vector(63 downto 0);
    input_1_input_count           : in std_logic_vector(3 downto 0);
    input_1_input_unl_valid       : in std_logic;
    input_1_input_unl_ready       : out std_logic;
    input_1_input_unl_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    input_1_input_cmd_valid       : out std_logic;
    input_1_input_cmd_ready       : in std_logic;
    input_1_input_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_1_input_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_1_input_cmd_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    input_2_input_valid           : in std_logic;
    input_2_input_ready           : out std_logic;
    input_2_input_dvalid          : in std_logic;
    input_2_input_last            : in std_logic;
    input_2_input                 : in std_logic_vector(63 downto 0);
    input_2_input_count           : in std_logic_vector(3 downto 0);
    input_2_input_unl_valid       : in std_logic;
    input_2_input_unl_ready       : out std_logic;
    input_2_input_unl_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    input_2_input_cmd_valid       : out std_logic;
    input_2_input_cmd_ready       : in std_logic;
    input_2_input_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_2_input_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    input_2_input_cmd_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_1_voltage_valid        : out std_logic;
    output_1_voltage_ready        : in std_logic;
    output_1_voltage_dvalid       : out std_logic;
    output_1_voltage_last         : out std_logic;
    output_1_voltage_length       : out std_logic_vector(31 downto 0);
    output_1_voltage_count        : out std_logic_vector(0 downto 0);
    output_1_voltage_item_valid   : out std_logic;
    output_1_voltage_item_ready   : in std_logic;
    output_1_voltage_item_dvalid  : out std_logic;
    output_1_voltage_item_last    : out std_logic;
    output_1_voltage_item         : out std_logic_vector(63 downto 0);
    output_1_voltage_item_count   : out std_logic_vector(0 downto 0);
    output_1_voltage_unl_valid    : in std_logic;
    output_1_voltage_unl_ready    : out std_logic;
    output_1_voltage_unl_tag      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_1_voltage_cmd_valid    : out std_logic;
    output_1_voltage_cmd_ready    : in std_logic;
    output_1_voltage_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_1_voltage_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_1_voltage_cmd_tag      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_2_voltage_valid        : out std_logic;
    output_2_voltage_ready        : in std_logic;
    output_2_voltage_dvalid       : out std_logic;
    output_2_voltage_last         : out std_logic;
    output_2_voltage_length       : out std_logic_vector(31 downto 0);
    output_2_voltage_count        : out std_logic_vector(0 downto 0);
    output_2_voltage_item_valid   : out std_logic;
    output_2_voltage_item_ready   : in std_logic;
    output_2_voltage_item_dvalid  : out std_logic;
    output_2_voltage_item_last    : out std_logic;
    output_2_voltage_item         : out std_logic_vector(63 downto 0);
    output_2_voltage_item_count   : out std_logic_vector(0 downto 0);
    output_2_voltage_unl_valid    : in std_logic;
    output_2_voltage_unl_ready    : out std_logic;
    output_2_voltage_unl_tag      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    output_2_voltage_cmd_valid    : out std_logic;
    output_2_voltage_cmd_ready    : in std_logic;
    output_2_voltage_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_2_voltage_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
    output_2_voltage_cmd_tag      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    start                         : in std_logic;
    stop                          : in std_logic;
    reset                         : in std_logic;
    idle                          : out std_logic;
    busy                          : out std_logic;
    done                          : out std_logic;
    result                        : out std_logic_vector(63 downto 0);
    input_1_firstidx              : in std_logic_vector(31 downto 0);
    input_1_lastidx               : in std_logic_vector(31 downto 0);
    input_2_firstidx              : in std_logic_vector(31 downto 0);
    input_2_lastidx               : in std_logic_vector(31 downto 0);
    output_1_firstidx             : in std_logic_vector(31 downto 0);
    output_1_lastidx              : in std_logic_vector(31 downto 0);
    output_2_firstidx             : in std_logic_vector(31 downto 0);
    output_2_lastidx              : in std_logic_vector(31 downto 0);
    ext_platform_complete_req     : out std_logic;
    ext_platform_complete_ack     : in std_logic
  );
end entity;

architecture Implementation of battery_status_2 is

  -- elements per cycle of input stream
  -- matches the value set in the schema (generate.py)
  constant EPC : natural := 8;

  type state_t is (
    STATE_IDLE,           -- idle
    STATE_REQ_READ_1,     -- send read request
    STATE_REQ_WRITE_1,    -- send write request
    STATE_REQ_READ_2,     -- send read request
    STATE_REQ_WRITE_2,    -- send write request
    STATE_UNLOCK_READ_1,  -- unlock read
    STATE_UNLOCK_READ_2,  -- unlock read
    STATE_UNLOCK_WRITE_1, -- unlock write
    STATE_UNLOCK_WRITE_2, -- unlock write
    STATE_FENCE,          -- write fence
    STATE_DONE            -- done
  );

  -- state signals
  signal state, state_next                                : state_t;

  -- parser output signals
  signal json_out_valid_1, json_out_valid_2               : std_logic;
  signal json_out_ready_1, json_out_ready_2               : std_logic;
  signal json_out_data_1, json_out_data_2                 : std_logic_vector(63 downto 0);
  signal json_out_last_1, json_out_last_2                 : std_logic_vector(2 downto 0);
  signal json_out_strb_1, json_out_strb_2                 : std_logic;

  signal int_input_input_ready_1, int_input_input_ready_2 : std_logic;

  signal strb_1, strb_2                                   : std_logic_vector(EPC - 1 downto 0);
  signal int_in_last_1, int_in_last_2                     : std_logic_vector(2 * EPC - 1 downto 0);

  signal cmd_complete_1, cmd_complete_2                   : std_logic;

  signal record_counter_1, record_counter_2               : unsigned(31 downto 0);

begin

  counter_1 : process (kcd_clk)
    is
  begin
    if rising_edge(kcd_clk) then
      if json_out_ready_1 = '1' and json_out_valid_1 = '1' and json_out_last_1(1) = '1' then
        record_counter_1 <= record_counter_1 + 1;
      end if;
      if kcd_reset = '1' or reset = '1' then
        record_counter_1 <= (others => '0');
      end if;
    end if;
  end process;

  counter_2 : process (kcd_clk)
    is
  begin
    if rising_edge(kcd_clk) then
      if json_out_ready_2 = '1' and json_out_valid_2 = '1' and json_out_last_2(1) = '1' then
        record_counter_2 <= record_counter_2 + 1;
      end if;
      if kcd_reset = '1' or reset = '1' then
        record_counter_2 <= (others => '0');
      end if;
    end if;
  end process;

  result <= std_logic_vector(record_counter_2) & std_logic_vector(record_counter_1);

  comb : process (
    start,
    reset,
    state,
    input_1_firstidx,
    input_1_lastidx,
    output_1_firstidx,
    output_1_lastidx,
    int_input_input_ready_1,
    input_1_input_cmd_ready,
    output_1_voltage_cmd_ready,
    input_1_input_unl_valid,
    output_1_voltage_unl_valid,
    input_2_firstidx,
    input_2_lastidx,
    output_2_firstidx,
    output_2_lastidx,
    int_input_input_ready_2,
    input_2_input_cmd_ready,
    output_2_voltage_cmd_ready,
    input_2_input_unl_valid,
    output_2_voltage_unl_valid,
    ext_platform_complete_ack
    ) is
  begin

    -- read request defaults
    input_1_input_cmd_valid       <= '0';
    input_1_input_cmd_firstIdx    <= input_1_firstidx;
    input_1_input_cmd_lastIdx     <= input_1_lastidx;
    input_1_input_cmd_tag         <= (others => '0');
    input_1_input_unl_ready       <= '0';

    input_2_input_cmd_valid       <= '0';
    input_2_input_cmd_firstIdx    <= input_2_firstidx;
    input_2_input_cmd_lastIdx     <= input_2_lastidx;
    input_2_input_cmd_tag         <= (others => '0');
    input_2_input_unl_ready       <= '0';

    -- write request defaults
    output_1_voltage_cmd_valid    <= '0';
    output_1_voltage_cmd_firstIdx <= output_1_firstidx;
    output_1_voltage_cmd_lastIdx  <= output_1_lastidx;
    output_1_voltage_cmd_tag      <= (others => '0');
    output_1_voltage_unl_ready    <= '0';

    output_2_voltage_cmd_valid    <= '0';
    output_2_voltage_cmd_firstIdx <= output_2_firstidx;
    output_2_voltage_cmd_lastIdx  <= output_2_lastidx;
    output_2_voltage_cmd_tag      <= (others => '0');
    output_2_voltage_unl_ready    <= '0';

    -- next state is the same if not changed
    state_next                    <= state;

    -- internal signal
    input_1_input_ready           <= int_input_input_ready_1;
    input_2_input_ready           <= int_input_input_ready_2;

    ext_platform_complete_req     <= '0';

    case state is

        -- wait for start signal
      when STATE_IDLE =>
        done <= '0';
        busy <= '0';
        idle <= '1';

        if start = '1' then
          state_next <= STATE_REQ_READ_1;
        end if;

        -- send read request
      when STATE_REQ_READ_1 =>
        done                    <= '0';
        busy                    <= '1';
        idle                    <= '0';

        input_1_input_cmd_valid <= '1';

        -- handshake
        if input_1_input_cmd_ready = '1' then
          state_next <= STATE_REQ_READ_2;
        end if;

        -- send read request
      when STATE_REQ_READ_2 =>
        done                    <= '0';
        busy                    <= '1';
        idle                    <= '0';

        input_2_input_cmd_valid <= '1';

        -- handshake
        if input_2_input_cmd_ready = '1' then
          state_next <= STATE_REQ_WRITE_1;
        end if;

        -- send write request
      when STATE_REQ_WRITE_1 =>
        done                       <= '0';
        busy                       <= '1';
        idle                       <= '0';

        output_1_voltage_cmd_valid <= '1';

        -- handshake
        if output_1_voltage_cmd_ready = '1' then
          state_next <= STATE_REQ_WRITE_2;
          -- state_next <= STATE_UNLOCK_READ;
        end if;

        -- send write request
      when STATE_REQ_WRITE_2 =>
        done                       <= '0';
        busy                       <= '1';
        idle                       <= '0';

        output_2_voltage_cmd_valid <= '1';

        -- handshake
        if output_2_voltage_cmd_ready = '1' then
          state_next <= STATE_UNLOCK_READ_1;
        end if;

        -- unlock read
      when STATE_UNLOCK_READ_1 =>
        done <= '0';
        busy <= '1';
        idle <= '0';

        if input_1_input_unl_valid = '1' then
          input_1_input_unl_ready <= '1';
          state_next              <= STATE_UNLOCK_READ_2;
          -- state_next            <= STATE_UNLOCK_WRITE;
        end if;

        -- unlock read
      when STATE_UNLOCK_READ_2 =>
        done <= '0';
        busy <= '1';
        idle <= '0';

        if input_2_input_unl_valid = '1' then
          input_2_input_unl_ready <= '1';
          state_next              <= STATE_UNLOCK_WRITE_1;
        end if;

        -- unlock write
      when STATE_UNLOCK_WRITE_1 =>
        done <= '0';
        busy <= '1';
        idle <= '0';

        if output_1_voltage_unl_valid = '1' then
          output_1_voltage_unl_ready <= '1';
          state_next                 <= STATE_UNLOCK_WRITE_2;
          -- state_next               <= STATE_FENCE;
        end if;

        -- unlock write
      when STATE_UNLOCK_WRITE_2 =>
        done <= '0';
        busy <= '1';
        idle <= '0';

        if output_2_voltage_unl_valid = '1' then
          output_2_voltage_unl_ready <= '1';
          state_next                 <= STATE_FENCE;
        end if;

      when STATE_FENCE =>
        done                      <= '0';
        busy                      <= '1';
        idle                      <= '0';

        ext_platform_complete_req <= '1';
        if ext_platform_complete_ack = '1' then
          state_next <= STATE_DONE;
        end if;

        -- wait for kernel reset
      when STATE_DONE =>
        done <= '1';
        busy <= '0';
        idle <= '1';

        if reset = '1' then
          state_next <= STATE_IDLE;
        end if;

    end case;

  end process;

  seq : process (kcd_clk)
  begin
    if rising_edge(kcd_clk) then
      state <= state_next;

      if kcd_reset = '1' then
        state <= STATE_IDLE;
      end if;

    end if;
  end process;

  tydi_strb : process (input_1_input_dvalid, input_1_input_count, input_2_input_dvalid, input_2_input_count)
  begin
    strb_1 <= (others => '0');
    strb_2 <= (others => '0');
    for i in strb_1'range loop
      if unsigned(input_1_input_count) = 0 or i < unsigned(input_1_input_count) then
        strb_1(i) <= input_1_input_dvalid;
      end if;
    end loop;
    for i in strb_2'range loop
      if unsigned(input_2_input_count) = 0 or i < unsigned(input_2_input_count) then
        strb_2(i) <= input_2_input_dvalid;
      end if;
    end loop;
  end process;

  int_in_last_proc : process (input_1_input_last, input_2_input_last)
  begin
    int_in_last_1              <= (others => '0');
    -- all records are currently sent in one transfer, so there's no difference
    -- between the two dimensions going into the parser.
    int_in_last_1(EPC * 2 - 2) <= input_1_input_last;
    int_in_last_1(EPC * 2 - 1) <= input_1_input_last;

    int_in_last_2              <= (others => '0');
    -- all records are currently sent in one transfer, so there's no difference
    -- between the two dimensions going into the parser.
    int_in_last_2(EPC * 2 - 2) <= input_2_input_last;
    int_in_last_2(EPC * 2 - 1) <= input_2_input_last;
  end process;

  battery_status_parser_1 : BattSchemaParser
  generic map(
    EPC                   => EPC,
    INT_WIDTH             => 64,
    INT_P_PIPELINE_STAGES => 4,
    END_REQ_EN            => false
  )
  port map(
    clk       => kcd_clk,
    reset     => kcd_reset,
    in_valid  => input_1_input_valid,
    in_ready  => int_input_input_ready_1,
    in_data   => input_1_input,
    in_last   => int_in_last_1,
    in_stai => (others => '0'),
    in_endi => (others => '1'),
    in_strb   => strb_1,
    end_req   => '0',  -- not implemented
    end_ack   => open, -- not implemented
    out_valid => json_out_valid_1,
    out_ready => json_out_ready_1,
    out_data  => json_out_data_1,
    out_last  => json_out_last_1,
    out_strb  => json_out_strb_1
  );
  battery_status_parser_2 : BattSchemaParser
  generic map(
    EPC                   => EPC,
    INT_WIDTH             => 64,
    INT_P_PIPELINE_STAGES => 4,
    END_REQ_EN            => false
  )
  port map(
    clk       => kcd_clk,
    reset     => kcd_reset,
    in_valid  => input_2_input_valid,
    in_ready  => int_input_input_ready_2,
    in_data   => input_2_input,
    in_last   => int_in_last_2,
    in_stai => (others => '0'),
    in_endi => (others => '1'),
    in_strb   => strb_2,
    end_req   => '0',  -- not implemented
    end_ack   => open, -- not implemented
    out_valid => json_out_valid_2,
    out_ready => json_out_ready_2,
    out_data  => json_out_data_2,
    out_last  => json_out_last_2,
    out_strb  => json_out_strb_2
  );

  convert_proc : process (kcd_clk) is

    type input_holding_reg_type is record
      valid         : std_logic;
      dvalid        : std_logic;
      data          : std_logic_vector(63 downto 0);
      end_of_array  : std_logic;
      end_of_object : std_logic;
      end_of_query  : std_logic;
    end record;
    variable i1, i2 : input_holding_reg_type;

    type count_output_holding_reg_type is record
      valid  : std_logic;
      dvalid : std_logic;
      data   : std_logic_vector(31 downto 0);
      last   : std_logic;
    end record;
    variable oc1, oc2 : count_output_holding_reg_type;

    type element_output_holding_reg_type is record
      valid  : std_logic;
      dvalid : std_logic;
      data   : std_logic_vector(63 downto 0);
      last   : std_logic;
    end record;
    variable oe1, oe2       : element_output_holding_reg_type;

    -- Current element count for length stream.
    variable count1, count2 : unsigned(31 downto 0) := (others => '0');

  begin

    if rising_edge(kcd_clk) then
      cmd_complete_1 <= '0';
      cmd_complete_2 <= '0';

      if i1.valid = '0' then
        i1.valid         := json_out_valid_1;
        i1.dvalid        := json_out_strb_1;
        i1.data          := json_out_data_1;
        i1.end_of_array  := json_out_last_1(0);
        i1.end_of_object := json_out_last_1(1);
        i1.end_of_query  := json_out_last_1(2);
      end if;

      if i2.valid = '0' then
        i2.valid         := json_out_valid_2;
        i2.dvalid        := json_out_strb_2;
        i2.data          := json_out_data_2;
        i2.end_of_array  := json_out_last_2(0);
        i2.end_of_object := json_out_last_2(1);
        i2.end_of_query  := json_out_last_2(2);
      end if;

      if output_1_voltage_ready = '1' then
        oc1.valid := '0';
      end if;
      if output_2_voltage_ready = '1' then
        oc2.valid := '0';
      end if;

      if output_1_voltage_item_ready = '1' then
        oe1.valid := '0';
      end if;
      if output_2_voltage_item_ready = '1' then
        oe2.valid := '0';
      end if;

      if i1.valid = '1' and oc1.valid = '0' and oe1.valid = '0' then
        oe1.dvalid := '0';
        oe1.last   := '0';
        oc1.dvalid := '0';
        oc1.last   := '0';

        -- If the data is valid, forward it and increment the element counter.
        if i1.dvalid = '1' then
          -- oe.valid  := '1';
          oe1.dvalid := '1';
          oe1.data   := i1.data;
          count1     := count1 + 1;
        end if;

        -- If this is the end of the current JSON object, send last to the
        -- element stream and send the element count to the length stream.
        -- We could also use end_of_array here; for valid JSON these should be
        -- equivalent.
        if i1.end_of_object = '1' then
          -- oc.valid  := '1';
          oc1.dvalid := '1';
          oc1.data   := std_logic_vector(count1);
          count1     := (others => '0');
        end if;

        -- If this is the end of the current command, send last to the length
        -- stream, and send a strobe to the state machine that indicates
        -- completion.
        if i1.end_of_query = '1' then
          -- oe.valid := '1';
          oe1.last := '1';
          -- oc.valid := '1';
          oc1.last := '1';
          cmd_complete_1 <= '0';
        end if;

        oe1.valid := i1.dvalid or i1.end_of_query;
        oc1.valid := i1.end_of_object or i1.end_of_query;

        -- clear holding register
        i1.valid  := '0';

      end if;

      if kcd_reset = '1' then
        i1.valid  := '0';
        oc1.valid := '0';
        oe1.valid := '0';
        count1    := (others => '0');
        cmd_complete_1 <= '0';
      end if;

      json_out_ready_1             <= not i1.valid;

      output_1_voltage_valid       <= oc1.valid;
      output_1_voltage_dvalid      <= oc1.dvalid;
      output_1_voltage_last        <= oc1.last;
      output_1_voltage_length      <= oc1.data;
      output_1_voltage_count       <= "1";

      output_1_voltage_item_valid  <= oe1.valid;
      output_1_voltage_item_dvalid <= oe1.dvalid;
      output_1_voltage_item_last   <= oe1.last;
      output_1_voltage_item        <= oe1.data;
      output_1_voltage_item_count  <= "1";

      if i2.valid = '1' and oc2.valid = '0' and oe2.valid = '0' then
        oe2.dvalid := '0';
        oe2.last   := '0';
        oc2.dvalid := '0';
        oc2.last   := '0';

        -- If the data is valid, forward it and increment the element counter.
        if i2.dvalid = '1' then
          -- oe.valid  := '1';
          oe2.dvalid := '1';
          oe2.data   := i2.data;
          count2     := count2 + 1;
        end if;

        -- If this is the end of the current JSON object, send last to the
        -- element stream and send the element count to the length stream.
        -- We could also use end_of_array here; for valid JSON these should be
        -- equivalent.
        if i2.end_of_object = '1' then
          -- oc.valid  := '1';
          oc2.dvalid := '1';
          oc2.data   := std_logic_vector(count2);
          count2     := (others => '0');
        end if;

        -- If this is the end of the current command, send last to the length
        -- stream, and send a strobe to the state machine that indicates
        -- completion.
        if i2.end_of_query = '1' then
          -- oe.valid := '1';
          oe2.last := '1';
          -- oc.valid := '1';
          oc2.last := '1';
          cmd_complete_2 <= '0';
        end if;

        oe2.valid := i2.dvalid or i2.end_of_query;
        oc2.valid := i2.end_of_object or i2.end_of_query;

        -- clear holding register
        i2.valid  := '0';

      end if;

      if kcd_reset = '1' then
        i2.valid  := '0';
        oc2.valid := '0';
        oe2.valid := '0';
        count2    := (others => '0');
        cmd_complete_2 <= '0';
      end if;

      json_out_ready_2             <= not i2.valid;

      output_2_voltage_valid       <= oc2.valid;
      output_2_voltage_dvalid      <= oc2.dvalid;
      output_2_voltage_last        <= oc2.last;
      output_2_voltage_length      <= oc2.data;
      output_2_voltage_count       <= "1";

      output_2_voltage_item_valid  <= oe2.valid;
      output_2_voltage_item_dvalid <= oe2.dvalid;
      output_2_voltage_item_last   <= oe2.last;
      output_2_voltage_item        <= oe2.data;
      output_2_voltage_item_count  <= "1";

    end if;

  end process;

end architecture;